	mem(0) := To_stdlogicvector(X"0D");
	mem(1) := To_stdlogicvector(X"62");
	mem(2) := To_stdlogicvector(X"10");
	mem(3) := To_stdlogicvector(X"72");
	mem(4) := To_stdlogicvector(X"11");
	mem(5) := To_stdlogicvector(X"74");
	mem(6) := To_stdlogicvector(X"12");
	mem(7) := To_stdlogicvector(X"76");
	mem(8) := To_stdlogicvector(X"10");
	mem(9) := To_stdlogicvector(X"68");
	mem(10) := To_stdlogicvector(X"11");
	mem(11) := To_stdlogicvector(X"6A");
	mem(12) := To_stdlogicvector(X"12");
	mem(13) := To_stdlogicvector(X"6C");
	mem(14) := To_stdlogicvector(X"FF");
	mem(15) := To_stdlogicvector(X"0F");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"D0");
	mem(23) := To_stdlogicvector(X"BA");
	mem(24) := To_stdlogicvector(X"D1");
	mem(25) := To_stdlogicvector(X"BA");
	mem(26) := To_stdlogicvector(X"0D");
	mem(27) := To_stdlogicvector(X"60");
	mem(28) := To_stdlogicvector(X"D2");
	mem(29) := To_stdlogicvector(X"BA");
	mem(30) := To_stdlogicvector(X"D3");
	mem(31) := To_stdlogicvector(X"BA");
	mem(32) := To_stdlogicvector(X"D1");
	mem(33) := To_stdlogicvector(X"BA");
	mem(34) := To_stdlogicvector(X"D2");
	mem(35) := To_stdlogicvector(X"BA");
	mem(36) := To_stdlogicvector(X"D3");
	mem(37) := To_stdlogicvector(X"BA");
