	mem(0) := To_stdlogicvector(X"62");
	mem(1) := To_stdlogicvector(X"12");
	mem(2) := To_stdlogicvector(X"55");
	mem(3) := To_stdlogicvector(X"64");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"A1");
	mem(7) := To_stdlogicvector(X"16");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"00");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"E1");
	mem(21) := To_stdlogicvector(X"18");
	mem(22) := To_stdlogicvector(X"55");
	mem(23) := To_stdlogicvector(X"78");
	mem(24) := To_stdlogicvector(X"55");
	mem(25) := To_stdlogicvector(X"6A");
	mem(26) := To_stdlogicvector(X"00");
	mem(27) := To_stdlogicvector(X"00");
	mem(28) := To_stdlogicvector(X"00");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"00");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"00");
	mem(33) := To_stdlogicvector(X"00");
	mem(34) := To_stdlogicvector(X"00");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"55");
	mem(39) := To_stdlogicvector(X"6A");
	mem(40) := To_stdlogicvector(X"64");
	mem(41) := To_stdlogicvector(X"11");
	mem(42) := To_stdlogicvector(X"00");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"32");
	mem(45) := To_stdlogicvector(X"00");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"00");
	mem(49) := To_stdlogicvector(X"00");
	mem(50) := To_stdlogicvector(X"00");
	mem(51) := To_stdlogicvector(X"00");
	mem(52) := To_stdlogicvector(X"00");
	mem(53) := To_stdlogicvector(X"00");
	mem(54) := To_stdlogicvector(X"00");
	mem(55) := To_stdlogicvector(X"00");
	mem(56) := To_stdlogicvector(X"00");
	mem(57) := To_stdlogicvector(X"00");
