--
-- VHDL Architecture ece411.Memory.untitled
--
-- Created:
--          by - tkalbar2.stdt (eelnx13.ews.illinois.edu)
--          at - 23:22:59 09/01/10
--
-- using Mentor Graphics HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      ADDRESS   : IN     LC3b_word;
      DATAOUT   : IN     LC3b_word;
      MREAD_L   : IN     std_logic;
      MWRITEH_L : IN     std_logic;
      MWRITEL_L : IN     std_logic;
      RESET_L   : IN     std_logic;
      clk       : IN     std_logic;
      DATAIN    : OUT    LC3b_word;
      MRESP_H   : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - tkalbar2.ece411_G2 (eelnx34.ews.illinois.edu)
--          at - 23:54:29 10/19/10
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2005.3 (Build 75)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY ece411;

ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL PMADDRESS    : LC3b_word;
   SIGNAL PMREAD_L     : std_logic;
   SIGNAL PMWRITE_L    : std_logic;
   SIGNAL dirty        : std_logic;
   SIGNAL in_idlehit   : std_logic;
   SIGNAL in_load      : std_logic;
   SIGNAL in_writeback : std_logic;
   SIGNAL miss         : std_logic;
   SIGNAL pmdatain     : LC3b_oword;
   SIGNAL pmdataout    : LC3b_oword;
   SIGNAL pmresp_h     : std_logic;


   -- Component Declarations
   COMPONENT Cache_Controller
   PORT (
      RESET_L      : IN     std_logic ;
      clk          : IN     std_logic ;
      dirty        : IN     std_logic ;
      miss         : IN     std_logic ;
      pmresp_h     : IN     std_logic ;
      PMREAD_L     : OUT    std_logic ;
      PMWRITE_L    : OUT    std_logic ;
      in_idlehit   : OUT    std_logic ;
      in_load      : OUT    std_logic ;
      in_writeback : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Cache_Datapath
   PORT (
      ADDRESS      : IN     LC3b_word ;
      DATAOUT      : IN     LC3b_word ;
      MREAD_L      : IN     std_logic ;
      MWRITEH_L    : IN     std_logic ;
      MWRITEL_L    : IN     std_logic ;
      RESET_L      : IN     std_logic ;
      clk          : IN     std_logic ;
      in_idlehit   : IN     std_logic ;
      in_load      : IN     std_logic ;
      in_writeback : IN     std_logic ;
      pmdatain     : IN     LC3b_oword ;
      pmresp_h     : IN     std_logic ;
      DATAIN       : OUT    LC3b_word ;
      MRESP_H      : OUT    std_logic ;
      PMADDRESS    : OUT    LC3b_word ;
      dirty        : OUT    std_logic ;
      miss         : OUT    std_logic ;
      pmdataout    : OUT    LC3b_oword 
   );
   END COMPONENT;
   COMPONENT DRAMAuditor
   PORT (
      ADDRESS   : IN     LC3b_word ;
      MREAD_L   : IN     std_logic ;
      MWRITEH_L : IN     std_logic ;
      MWRITEL_L : IN     std_logic ;
      RESET_L   : IN     std_logic 
   );
   END COMPONENT;
   COMPONENT PDRAMAuditor
   PORT (
      PMADDRESS : IN     LC3b_word ;
      RESET_L   : IN     std_logic ;
      PMREAD_L  : IN     std_logic ;
      PMWRITE_L : IN     std_logic 
   );
   END COMPONENT;
   COMPONENT Physical_Memory
   PORT (
      PMADDRESS : IN     LC3b_word ;
      pmdataout : IN     LC3b_oword ;
      pmdatain  : OUT    LC3b_oword ;
      PMWRITE_L : IN     std_logic ;
      PMREAD_L  : IN     std_logic ;
      pmresp_h  : OUT    std_logic ;
      RESET_L   : IN     std_logic ;
      clk       : IN     std_logic 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Controller USE ENTITY ece411.Cache_Controller;
   FOR ALL : Cache_Datapath USE ENTITY ece411.Cache_Datapath;
   FOR ALL : DRAMAuditor USE ENTITY ece411.DRAMAuditor;
   FOR ALL : PDRAMAuditor USE ENTITY ece411.PDRAMAuditor;
   FOR ALL : Physical_Memory USE ENTITY ece411.Physical_Memory;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   Cache_Cont : Cache_Controller
      PORT MAP (
         RESET_L      => RESET_L,
         clk          => clk,
         dirty        => dirty,
         miss         => miss,
         pmresp_h     => pmresp_h,
         PMREAD_L     => PMREAD_L,
         PMWRITE_L    => PMWRITE_L,
         in_idlehit   => in_idlehit,
         in_load      => in_load,
         in_writeback => in_writeback
      );
   Cache_DP : Cache_Datapath
      PORT MAP (
         ADDRESS      => ADDRESS,
         DATAOUT      => DATAOUT,
         MREAD_L      => MREAD_L,
         MWRITEH_L    => MWRITEH_L,
         MWRITEL_L    => MWRITEL_L,
         RESET_L      => RESET_L,
         clk          => clk,
         in_idlehit   => in_idlehit,
         in_load      => in_load,
         in_writeback => in_writeback,
         pmdatain     => pmdatain,
         pmresp_h     => pmresp_h,
         DATAIN       => DATAIN,
         MRESP_H      => MRESP_H,
         PMADDRESS    => PMADDRESS,
         dirty        => dirty,
         miss         => miss,
         pmdataout    => pmdataout
      );
   U_1 : DRAMAuditor
      PORT MAP (
         ADDRESS   => ADDRESS,
         MREAD_L   => MREAD_L,
         MWRITEH_L => MWRITEH_L,
         MWRITEL_L => MWRITEL_L,
         RESET_L   => RESET_L
      );
   U_0 : PDRAMAuditor
      PORT MAP (
         PMADDRESS => PMADDRESS,
         RESET_L   => RESET_L,
         PMREAD_L  => PMREAD_L,
         PMWRITE_L => PMWRITE_L
      );
   PDRAM : Physical_Memory
      PORT MAP (
         PMADDRESS => PMADDRESS,
         pmdataout => pmdataout,
         pmdatain  => pmdatain,
         PMWRITE_L => PMWRITE_L,
         PMREAD_L  => PMREAD_L,
         pmresp_h  => pmresp_h,
         RESET_L   => RESET_L,
         clk       => clk
      );

END struct;
