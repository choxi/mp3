	mem(0) := To_stdlogicvector(X"7F");
	mem(1) := To_stdlogicvector(X"12");
	mem(2) := To_stdlogicvector(X"BF");
	mem(3) := To_stdlogicvector(X"14");
	mem(4) := To_stdlogicvector(X"14");
	mem(5) := To_stdlogicvector(X"2C");
	mem(6) := To_stdlogicvector(X"15");
	mem(7) := To_stdlogicvector(X"2E");
	mem(8) := To_stdlogicvector(X"14");
	mem(9) := To_stdlogicvector(X"22");
	mem(10) := To_stdlogicvector(X"15");
	mem(11) := To_stdlogicvector(X"24");
	mem(12) := To_stdlogicvector(X"16");
	mem(13) := To_stdlogicvector(X"3C");
	mem(14) := To_stdlogicvector(X"17");
	mem(15) := To_stdlogicvector(X"3E");
	mem(16) := To_stdlogicvector(X"0B");
	mem(17) := To_stdlogicvector(X"6A");
	mem(18) := To_stdlogicvector(X"FF");
	mem(19) := To_stdlogicvector(X"0F");
	mem(20) := To_stdlogicvector(X"0D");
	mem(21) := To_stdlogicvector(X"60");
	mem(22) := To_stdlogicvector(X"FF");
	mem(23) := To_stdlogicvector(X"FF");
