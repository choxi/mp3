	mem(0) := To_stdlogicvector(X"0B");
	mem(1) := To_stdlogicvector(X"62");
	mem(2) := To_stdlogicvector(X"0C");
	mem(3) := To_stdlogicvector(X"64");
	mem(4) := To_stdlogicvector(X"0D");
	mem(5) := To_stdlogicvector(X"66");
	mem(6) := To_stdlogicvector(X"40");
	mem(7) := To_stdlogicvector(X"68");
	mem(8) := To_stdlogicvector(X"80");
	mem(9) := To_stdlogicvector(X"6A");
	mem(10) := To_stdlogicvector(X"40");
	mem(11) := To_stdlogicvector(X"6C");
	mem(12) := To_stdlogicvector(X"C0");
	mem(13) := To_stdlogicvector(X"6E");
	mem(14) := To_stdlogicvector(X"40");
	mem(15) := To_stdlogicvector(X"60");
	mem(16) := To_stdlogicvector(X"C0");
	mem(17) := To_stdlogicvector(X"62");
	mem(18) := To_stdlogicvector(X"80");
	mem(19) := To_stdlogicvector(X"64");
	mem(20) := To_stdlogicvector(X"FF");
	mem(21) := To_stdlogicvector(X"0F");
	mem(22) := To_stdlogicvector(X"20");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"A0");
	mem(25) := To_stdlogicvector(X"00");
	mem(26) := To_stdlogicvector(X"20");
	mem(27) := To_stdlogicvector(X"01");
	mem(32) := To_stdlogicvector(X"11");
	mem(33) := To_stdlogicvector(X"11");
	mem(34) := To_stdlogicvector(X"00");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"00");
	mem(39) := To_stdlogicvector(X"00");
	mem(40) := To_stdlogicvector(X"00");
	mem(41) := To_stdlogicvector(X"00");
	mem(42) := To_stdlogicvector(X"00");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"00");
	mem(45) := To_stdlogicvector(X"00");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(160) := To_stdlogicvector(X"22");
	mem(161) := To_stdlogicvector(X"22");
	mem(162) := To_stdlogicvector(X"00");
	mem(163) := To_stdlogicvector(X"00");
	mem(164) := To_stdlogicvector(X"00");
	mem(165) := To_stdlogicvector(X"00");
	mem(166) := To_stdlogicvector(X"00");
	mem(167) := To_stdlogicvector(X"00");
	mem(168) := To_stdlogicvector(X"00");
	mem(169) := To_stdlogicvector(X"00");
	mem(170) := To_stdlogicvector(X"00");
	mem(171) := To_stdlogicvector(X"00");
	mem(172) := To_stdlogicvector(X"00");
	mem(173) := To_stdlogicvector(X"00");
	mem(174) := To_stdlogicvector(X"00");
	mem(175) := To_stdlogicvector(X"00");
	mem(288) := To_stdlogicvector(X"33");
	mem(289) := To_stdlogicvector(X"33");
	mem(290) := To_stdlogicvector(X"00");
	mem(291) := To_stdlogicvector(X"00");
	mem(292) := To_stdlogicvector(X"00");
	mem(293) := To_stdlogicvector(X"00");
	mem(294) := To_stdlogicvector(X"00");
	mem(295) := To_stdlogicvector(X"00");
	mem(296) := To_stdlogicvector(X"00");
	mem(297) := To_stdlogicvector(X"00");
	mem(298) := To_stdlogicvector(X"00");
	mem(299) := To_stdlogicvector(X"00");
	mem(300) := To_stdlogicvector(X"00");
	mem(301) := To_stdlogicvector(X"00");
	mem(302) := To_stdlogicvector(X"00");
	mem(303) := To_stdlogicvector(X"00");
