	mem(0) := To_stdlogicvector(X"00");
	mem(1) := To_stdlogicvector(X"00");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"06");
	mem(11) := To_stdlogicvector(X"E0");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"12");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"00");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"32");
	mem(25) := To_stdlogicvector(X"00");
	mem(26) := To_stdlogicvector(X"00");
	mem(27) := To_stdlogicvector(X"00");
	mem(28) := To_stdlogicvector(X"00");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"00");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"00");
	mem(33) := To_stdlogicvector(X"00");
	mem(34) := To_stdlogicvector(X"00");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"00");
