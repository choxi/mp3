	mem(0) := To_stdlogicvector(X"00");
	mem(1) := To_stdlogicvector(X"00");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"22");
	mem(7) := To_stdlogicvector(X"10");
	mem(8) := To_stdlogicvector(X"09");
	mem(9) := To_stdlogicvector(X"A2");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"00");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"FF");
	mem(17) := To_stdlogicvector(X"0F");
	mem(18) := To_stdlogicvector(X"DD");
	mem(19) := To_stdlogicvector(X"B4");
	mem(20) := To_stdlogicvector(X"1E");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"DD");
	mem(23) := To_stdlogicvector(X"B4");
	mem(24) := To_stdlogicvector(X"DD");
	mem(25) := To_stdlogicvector(X"B4");
	mem(26) := To_stdlogicvector(X"DD");
	mem(27) := To_stdlogicvector(X"B4");
	mem(28) := To_stdlogicvector(X"DD");
	mem(29) := To_stdlogicvector(X"B4");
	mem(30) := To_stdlogicvector(X"0D");
	mem(31) := To_stdlogicvector(X"60");
	mem(32) := To_stdlogicvector(X"DD");
	mem(33) := To_stdlogicvector(X"B4");
	mem(34) := To_stdlogicvector(X"DD");
	mem(35) := To_stdlogicvector(X"B4");
	mem(36) := To_stdlogicvector(X"DD");
	mem(37) := To_stdlogicvector(X"B4");
	mem(38) := To_stdlogicvector(X"DD");
	mem(39) := To_stdlogicvector(X"B4");
	mem(40) := To_stdlogicvector(X"DD");
	mem(41) := To_stdlogicvector(X"B4");
	mem(42) := To_stdlogicvector(X"DD");
	mem(43) := To_stdlogicvector(X"B4");
	mem(44) := To_stdlogicvector(X"DD");
	mem(45) := To_stdlogicvector(X"B4");
	mem(46) := To_stdlogicvector(X"DD");
	mem(47) := To_stdlogicvector(X"B4");
	mem(48) := To_stdlogicvector(X"DD");
	mem(49) := To_stdlogicvector(X"B4");
	mem(50) := To_stdlogicvector(X"DD");
	mem(51) := To_stdlogicvector(X"B4");
	mem(52) := To_stdlogicvector(X"DD");
	mem(53) := To_stdlogicvector(X"B4");
	mem(54) := To_stdlogicvector(X"DD");
	mem(55) := To_stdlogicvector(X"B4");
