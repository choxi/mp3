	mem(0) := To_stdlogicvector(X"2F");
	mem(1) := To_stdlogicvector(X"E0");
	mem(2) := To_stdlogicvector(X"6E");
	mem(3) := To_stdlogicvector(X"E2");
	mem(4) := To_stdlogicvector(X"AD");
	mem(5) := To_stdlogicvector(X"E4");
	mem(6) := To_stdlogicvector(X"8A");
	mem(7) := To_stdlogicvector(X"6E");
	mem(8) := To_stdlogicvector(X"4B");
	mem(9) := To_stdlogicvector(X"6E");
	mem(10) := To_stdlogicvector(X"88");
	mem(11) := To_stdlogicvector(X"6C");
	mem(12) := To_stdlogicvector(X"0E");
	mem(13) := To_stdlogicvector(X"6E");
	mem(14) := To_stdlogicvector(X"0E");
	mem(15) := To_stdlogicvector(X"6C");
	mem(16) := To_stdlogicvector(X"4F");
	mem(17) := To_stdlogicvector(X"6C");
	mem(18) := To_stdlogicvector(X"8C");
	mem(19) := To_stdlogicvector(X"6C");
	mem(20) := To_stdlogicvector(X"8C");
	mem(21) := To_stdlogicvector(X"6C");
	mem(22) := To_stdlogicvector(X"8C");
	mem(23) := To_stdlogicvector(X"6C");
	mem(24) := To_stdlogicvector(X"81");
	mem(25) := To_stdlogicvector(X"6A");
	mem(26) := To_stdlogicvector(X"46");
	mem(27) := To_stdlogicvector(X"28");
	mem(28) := To_stdlogicvector(X"44");
	mem(29) := To_stdlogicvector(X"78");
	mem(30) := To_stdlogicvector(X"83");
	mem(31) := To_stdlogicvector(X"6A");
	mem(32) := To_stdlogicvector(X"4A");
	mem(33) := To_stdlogicvector(X"32");
	mem(34) := To_stdlogicvector(X"42");
	mem(35) := To_stdlogicvector(X"72");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"34");
	mem(38) := To_stdlogicvector(X"61");
	mem(39) := To_stdlogicvector(X"18");
	mem(40) := To_stdlogicvector(X"0A");
	mem(41) := To_stdlogicvector(X"39");
	mem(42) := To_stdlogicvector(X"02");
	mem(43) := To_stdlogicvector(X"E0");
	mem(44) := To_stdlogicvector(X"29");
	mem(45) := To_stdlogicvector(X"0E");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"0D");
	mem(49) := To_stdlogicvector(X"60");
	mem(50) := To_stdlogicvector(X"0D");
	mem(51) := To_stdlogicvector(X"60");
	mem(52) := To_stdlogicvector(X"0D");
	mem(53) := To_stdlogicvector(X"60");
	mem(54) := To_stdlogicvector(X"0D");
	mem(55) := To_stdlogicvector(X"60");
	mem(56) := To_stdlogicvector(X"0D");
	mem(57) := To_stdlogicvector(X"60");
	mem(58) := To_stdlogicvector(X"0D");
	mem(59) := To_stdlogicvector(X"60");
	mem(60) := To_stdlogicvector(X"0D");
	mem(61) := To_stdlogicvector(X"60");
	mem(62) := To_stdlogicvector(X"0D");
	mem(63) := To_stdlogicvector(X"60");
	mem(64) := To_stdlogicvector(X"C2");
	mem(65) := To_stdlogicvector(X"00");
	mem(66) := To_stdlogicvector(X"48");
	mem(67) := To_stdlogicvector(X"01");
	mem(68) := To_stdlogicvector(X"22");
	mem(69) := To_stdlogicvector(X"11");
	mem(70) := To_stdlogicvector(X"44");
	mem(71) := To_stdlogicvector(X"33");
	mem(72) := To_stdlogicvector(X"66");
	mem(73) := To_stdlogicvector(X"55");
	mem(74) := To_stdlogicvector(X"88");
	mem(75) := To_stdlogicvector(X"77");
	mem(76) := To_stdlogicvector(X"AA");
	mem(77) := To_stdlogicvector(X"99");
	mem(78) := To_stdlogicvector(X"CC");
	mem(79) := To_stdlogicvector(X"BB");
	mem(80) := To_stdlogicvector(X"0D");
	mem(81) := To_stdlogicvector(X"60");
	mem(82) := To_stdlogicvector(X"0D");
	mem(83) := To_stdlogicvector(X"60");
	mem(84) := To_stdlogicvector(X"0D");
	mem(85) := To_stdlogicvector(X"60");
	mem(86) := To_stdlogicvector(X"0D");
	mem(87) := To_stdlogicvector(X"60");
	mem(88) := To_stdlogicvector(X"0D");
	mem(89) := To_stdlogicvector(X"60");
	mem(90) := To_stdlogicvector(X"0D");
	mem(91) := To_stdlogicvector(X"60");
	mem(92) := To_stdlogicvector(X"0D");
	mem(93) := To_stdlogicvector(X"60");
	mem(94) := To_stdlogicvector(X"0D");
	mem(95) := To_stdlogicvector(X"60");
	mem(96) := To_stdlogicvector(X"6D");
	mem(97) := To_stdlogicvector(X"66");
	mem(98) := To_stdlogicvector(X"7D");
	mem(99) := To_stdlogicvector(X"67");
	mem(100) := To_stdlogicvector(X"8D");
	mem(101) := To_stdlogicvector(X"68");
	mem(102) := To_stdlogicvector(X"9D");
	mem(103) := To_stdlogicvector(X"69");
	mem(104) := To_stdlogicvector(X"AD");
	mem(105) := To_stdlogicvector(X"6A");
	mem(106) := To_stdlogicvector(X"BD");
	mem(107) := To_stdlogicvector(X"6B");
	mem(108) := To_stdlogicvector(X"CD");
	mem(109) := To_stdlogicvector(X"6C");
	mem(110) := To_stdlogicvector(X"DD");
	mem(111) := To_stdlogicvector(X"6D");
	mem(112) := To_stdlogicvector(X"0D");
	mem(113) := To_stdlogicvector(X"60");
	mem(114) := To_stdlogicvector(X"0D");
	mem(115) := To_stdlogicvector(X"60");
	mem(116) := To_stdlogicvector(X"0D");
	mem(117) := To_stdlogicvector(X"60");
	mem(118) := To_stdlogicvector(X"0D");
	mem(119) := To_stdlogicvector(X"60");
	mem(120) := To_stdlogicvector(X"0D");
	mem(121) := To_stdlogicvector(X"60");
	mem(122) := To_stdlogicvector(X"0D");
	mem(123) := To_stdlogicvector(X"60");
	mem(124) := To_stdlogicvector(X"0D");
	mem(125) := To_stdlogicvector(X"60");
	mem(126) := To_stdlogicvector(X"0D");
	mem(127) := To_stdlogicvector(X"60");
	mem(128) := To_stdlogicvector(X"17");
	mem(129) := To_stdlogicvector(X"E2");
	mem(130) := To_stdlogicvector(X"56");
	mem(131) := To_stdlogicvector(X"E4");
	mem(132) := To_stdlogicvector(X"10");
	mem(133) := To_stdlogicvector(X"70");
	mem(134) := To_stdlogicvector(X"51");
	mem(135) := To_stdlogicvector(X"72");
	mem(136) := To_stdlogicvector(X"92");
	mem(137) := To_stdlogicvector(X"74");
	mem(138) := To_stdlogicvector(X"14");
	mem(139) := To_stdlogicvector(X"74");
	mem(140) := To_stdlogicvector(X"51");
	mem(141) := To_stdlogicvector(X"6E");
	mem(142) := To_stdlogicvector(X"95");
	mem(143) := To_stdlogicvector(X"6A");
	mem(144) := To_stdlogicvector(X"12");
	mem(145) := To_stdlogicvector(X"6C");
	mem(146) := To_stdlogicvector(X"56");
	mem(147) := To_stdlogicvector(X"2A");
	mem(148) := To_stdlogicvector(X"A1");
	mem(149) := To_stdlogicvector(X"18");
	mem(150) := To_stdlogicvector(X"12");
	mem(151) := To_stdlogicvector(X"2D");
	mem(152) := To_stdlogicvector(X"46");
	mem(153) := To_stdlogicvector(X"1D");
	mem(154) := To_stdlogicvector(X"08");
	mem(155) := To_stdlogicvector(X"AA");
	mem(156) := To_stdlogicvector(X"46");
	mem(157) := To_stdlogicvector(X"1D");
	mem(158) := To_stdlogicvector(X"09");
	mem(159) := To_stdlogicvector(X"BC");
	mem(160) := To_stdlogicvector(X"E0");
	mem(161) := To_stdlogicvector(X"56");
	mem(162) := To_stdlogicvector(X"ED");
	mem(163) := To_stdlogicvector(X"16");
	mem(164) := To_stdlogicvector(X"00");
	mem(165) := To_stdlogicvector(X"3C");
	mem(166) := To_stdlogicvector(X"21");
	mem(167) := To_stdlogicvector(X"18");
	mem(168) := To_stdlogicvector(X"00");
	mem(169) := To_stdlogicvector(X"29");
	mem(170) := To_stdlogicvector(X"05");
	mem(171) := To_stdlogicvector(X"78");
	mem(172) := To_stdlogicvector(X"29");
	mem(173) := To_stdlogicvector(X"0E");
	mem(174) := To_stdlogicvector(X"00");
	mem(175) := To_stdlogicvector(X"00");
	mem(176) := To_stdlogicvector(X"20");
	mem(177) := To_stdlogicvector(X"52");
	mem(178) := To_stdlogicvector(X"20");
	mem(179) := To_stdlogicvector(X"52");
	mem(180) := To_stdlogicvector(X"20");
	mem(181) := To_stdlogicvector(X"52");
	mem(182) := To_stdlogicvector(X"20");
	mem(183) := To_stdlogicvector(X"52");
	mem(184) := To_stdlogicvector(X"20");
	mem(185) := To_stdlogicvector(X"52");
	mem(186) := To_stdlogicvector(X"20");
	mem(187) := To_stdlogicvector(X"52");
	mem(188) := To_stdlogicvector(X"20");
	mem(189) := To_stdlogicvector(X"52");
	mem(190) := To_stdlogicvector(X"20");
	mem(191) := To_stdlogicvector(X"52");
	mem(192) := To_stdlogicvector(X"20");
	mem(193) := To_stdlogicvector(X"52");
	mem(194) := To_stdlogicvector(X"20");
	mem(195) := To_stdlogicvector(X"52");
	mem(196) := To_stdlogicvector(X"20");
	mem(197) := To_stdlogicvector(X"52");
	mem(198) := To_stdlogicvector(X"20");
	mem(199) := To_stdlogicvector(X"52");
	mem(200) := To_stdlogicvector(X"20");
	mem(201) := To_stdlogicvector(X"52");
	mem(202) := To_stdlogicvector(X"20");
	mem(203) := To_stdlogicvector(X"52");
	mem(204) := To_stdlogicvector(X"20");
	mem(205) := To_stdlogicvector(X"52");
	mem(206) := To_stdlogicvector(X"20");
	mem(207) := To_stdlogicvector(X"52");
	mem(208) := To_stdlogicvector(X"20");
	mem(209) := To_stdlogicvector(X"52");
	mem(210) := To_stdlogicvector(X"20");
	mem(211) := To_stdlogicvector(X"52");
	mem(212) := To_stdlogicvector(X"20");
	mem(213) := To_stdlogicvector(X"52");
	mem(214) := To_stdlogicvector(X"20");
	mem(215) := To_stdlogicvector(X"52");
	mem(216) := To_stdlogicvector(X"20");
	mem(217) := To_stdlogicvector(X"52");
	mem(218) := To_stdlogicvector(X"20");
	mem(219) := To_stdlogicvector(X"52");
	mem(220) := To_stdlogicvector(X"20");
	mem(221) := To_stdlogicvector(X"52");
	mem(222) := To_stdlogicvector(X"20");
	mem(223) := To_stdlogicvector(X"52");
	mem(224) := To_stdlogicvector(X"A0");
	mem(225) := To_stdlogicvector(X"5A");
	mem(226) := To_stdlogicvector(X"B0");
	mem(227) := To_stdlogicvector(X"5B");
	mem(228) := To_stdlogicvector(X"C0");
	mem(229) := To_stdlogicvector(X"5C");
	mem(230) := To_stdlogicvector(X"D0");
	mem(231) := To_stdlogicvector(X"5D");
	mem(232) := To_stdlogicvector(X"E0");
	mem(233) := To_stdlogicvector(X"5E");
	mem(234) := To_stdlogicvector(X"F0");
	mem(235) := To_stdlogicvector(X"5F");
	mem(236) := To_stdlogicvector(X"10");
	mem(237) := To_stdlogicvector(X"51");
	mem(238) := To_stdlogicvector(X"20");
	mem(239) := To_stdlogicvector(X"52");
	mem(240) := To_stdlogicvector(X"20");
	mem(241) := To_stdlogicvector(X"52");
	mem(242) := To_stdlogicvector(X"20");
	mem(243) := To_stdlogicvector(X"52");
	mem(244) := To_stdlogicvector(X"20");
	mem(245) := To_stdlogicvector(X"52");
	mem(246) := To_stdlogicvector(X"20");
	mem(247) := To_stdlogicvector(X"52");
	mem(248) := To_stdlogicvector(X"20");
	mem(249) := To_stdlogicvector(X"52");
	mem(250) := To_stdlogicvector(X"20");
	mem(251) := To_stdlogicvector(X"52");
	mem(252) := To_stdlogicvector(X"20");
	mem(253) := To_stdlogicvector(X"52");
	mem(254) := To_stdlogicvector(X"20");
	mem(255) := To_stdlogicvector(X"52");
	mem(256) := To_stdlogicvector(X"42");
	mem(257) := To_stdlogicvector(X"6A");
	mem(258) := To_stdlogicvector(X"01");
	mem(259) := To_stdlogicvector(X"68");
	mem(260) := To_stdlogicvector(X"00");
	mem(261) := To_stdlogicvector(X"6C");
	mem(262) := To_stdlogicvector(X"04");
	mem(263) := To_stdlogicvector(X"2C");
	mem(264) := To_stdlogicvector(X"86");
	mem(265) := To_stdlogicvector(X"68");
	mem(266) := To_stdlogicvector(X"FF");
	mem(267) := To_stdlogicvector(X"16");
	mem(268) := To_stdlogicvector(X"F9");
	mem(269) := To_stdlogicvector(X"03");
	mem(270) := To_stdlogicvector(X"FF");
	mem(271) := To_stdlogicvector(X"0F");
	mem(272) := To_stdlogicvector(X"DD");
	mem(273) := To_stdlogicvector(X"BA");
	mem(274) := To_stdlogicvector(X"DD");
	mem(275) := To_stdlogicvector(X"BA");
	mem(276) := To_stdlogicvector(X"2D");
	mem(277) := To_stdlogicvector(X"B2");
	mem(278) := To_stdlogicvector(X"3D");
	mem(279) := To_stdlogicvector(X"B3");
	mem(280) := To_stdlogicvector(X"4D");
	mem(281) := To_stdlogicvector(X"B4");
	mem(282) := To_stdlogicvector(X"5D");
	mem(283) := To_stdlogicvector(X"B5");
	mem(284) := To_stdlogicvector(X"6D");
	mem(285) := To_stdlogicvector(X"B6");
	mem(286) := To_stdlogicvector(X"7D");
	mem(287) := To_stdlogicvector(X"B7");
	mem(288) := To_stdlogicvector(X"8D");
	mem(289) := To_stdlogicvector(X"B8");
	mem(290) := To_stdlogicvector(X"9D");
	mem(291) := To_stdlogicvector(X"B9");
	mem(292) := To_stdlogicvector(X"AD");
	mem(293) := To_stdlogicvector(X"BA");
	mem(294) := To_stdlogicvector(X"BD");
	mem(295) := To_stdlogicvector(X"BB");
	mem(296) := To_stdlogicvector(X"CD");
	mem(297) := To_stdlogicvector(X"BC");
	mem(298) := To_stdlogicvector(X"DD");
	mem(299) := To_stdlogicvector(X"BD");
	mem(300) := To_stdlogicvector(X"ED");
	mem(301) := To_stdlogicvector(X"BE");
	mem(302) := To_stdlogicvector(X"FD");
	mem(303) := To_stdlogicvector(X"BF");
	mem(304) := To_stdlogicvector(X"AD");
	mem(305) := To_stdlogicvector(X"BA");
	mem(306) := To_stdlogicvector(X"AD");
	mem(307) := To_stdlogicvector(X"BA");
	mem(308) := To_stdlogicvector(X"AD");
	mem(309) := To_stdlogicvector(X"BA");
	mem(310) := To_stdlogicvector(X"AD");
	mem(311) := To_stdlogicvector(X"BA");
	mem(312) := To_stdlogicvector(X"AD");
	mem(313) := To_stdlogicvector(X"BA");
	mem(314) := To_stdlogicvector(X"AD");
	mem(315) := To_stdlogicvector(X"BA");
	mem(316) := To_stdlogicvector(X"AD");
	mem(317) := To_stdlogicvector(X"BA");
	mem(318) := To_stdlogicvector(X"AD");
	mem(319) := To_stdlogicvector(X"BA");
	mem(320) := To_stdlogicvector(X"AD");
	mem(321) := To_stdlogicvector(X"BA");
	mem(322) := To_stdlogicvector(X"AD");
	mem(323) := To_stdlogicvector(X"BA");
	mem(324) := To_stdlogicvector(X"AD");
	mem(325) := To_stdlogicvector(X"BA");
	mem(326) := To_stdlogicvector(X"AD");
	mem(327) := To_stdlogicvector(X"BA");
	mem(328) := To_stdlogicvector(X"AD");
	mem(329) := To_stdlogicvector(X"BA");
	mem(330) := To_stdlogicvector(X"AD");
	mem(331) := To_stdlogicvector(X"BA");
	mem(332) := To_stdlogicvector(X"AD");
	mem(333) := To_stdlogicvector(X"BA");
	mem(334) := To_stdlogicvector(X"AD");
	mem(335) := To_stdlogicvector(X"BA");
	mem(336) := To_stdlogicvector(X"AD");
	mem(337) := To_stdlogicvector(X"BA");
	mem(338) := To_stdlogicvector(X"AD");
	mem(339) := To_stdlogicvector(X"BA");
	mem(340) := To_stdlogicvector(X"AD");
	mem(341) := To_stdlogicvector(X"BA");
	mem(342) := To_stdlogicvector(X"AD");
	mem(343) := To_stdlogicvector(X"BA");
	mem(344) := To_stdlogicvector(X"AD");
	mem(345) := To_stdlogicvector(X"BA");
	mem(346) := To_stdlogicvector(X"AD");
	mem(347) := To_stdlogicvector(X"BA");
	mem(348) := To_stdlogicvector(X"AD");
	mem(349) := To_stdlogicvector(X"BA");
	mem(350) := To_stdlogicvector(X"AD");
	mem(351) := To_stdlogicvector(X"BA");
	mem(352) := To_stdlogicvector(X"8D");
	mem(353) := To_stdlogicvector(X"B8");
	mem(354) := To_stdlogicvector(X"9D");
	mem(355) := To_stdlogicvector(X"B9");
	mem(356) := To_stdlogicvector(X"AD");
	mem(357) := To_stdlogicvector(X"BA");
	mem(358) := To_stdlogicvector(X"BD");
	mem(359) := To_stdlogicvector(X"BB");
	mem(360) := To_stdlogicvector(X"CD");
	mem(361) := To_stdlogicvector(X"BC");
	mem(362) := To_stdlogicvector(X"DD");
	mem(363) := To_stdlogicvector(X"BD");
	mem(364) := To_stdlogicvector(X"ED");
	mem(365) := To_stdlogicvector(X"BE");
	mem(366) := To_stdlogicvector(X"FD");
	mem(367) := To_stdlogicvector(X"BF");
	mem(368) := To_stdlogicvector(X"DD");
	mem(369) := To_stdlogicvector(X"BA");
	mem(370) := To_stdlogicvector(X"DD");
	mem(371) := To_stdlogicvector(X"BA");
	mem(372) := To_stdlogicvector(X"DD");
	mem(373) := To_stdlogicvector(X"BA");
	mem(374) := To_stdlogicvector(X"DD");
	mem(375) := To_stdlogicvector(X"BA");
	mem(376) := To_stdlogicvector(X"DD");
	mem(377) := To_stdlogicvector(X"BA");
	mem(378) := To_stdlogicvector(X"DD");
	mem(379) := To_stdlogicvector(X"BA");
	mem(380) := To_stdlogicvector(X"DD");
	mem(381) := To_stdlogicvector(X"BA");
	mem(382) := To_stdlogicvector(X"DD");
	mem(383) := To_stdlogicvector(X"BA");
