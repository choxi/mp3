	mem(0) := To_stdlogicvector(X"1A");
	mem(1) := To_stdlogicvector(X"6A");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"1D");
	mem(13) := To_stdlogicvector(X"7A");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"00");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"1D");
	mem(25) := To_stdlogicvector(X"6C");
	mem(26) := To_stdlogicvector(X"00");
	mem(27) := To_stdlogicvector(X"00");
	mem(28) := To_stdlogicvector(X"00");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"00");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"00");
	mem(33) := To_stdlogicvector(X"00");
	mem(34) := To_stdlogicvector(X"00");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"F9");
	mem(39) := To_stdlogicvector(X"0F");
	mem(40) := To_stdlogicvector(X"00");
	mem(41) := To_stdlogicvector(X"00");
	mem(42) := To_stdlogicvector(X"00");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"00");
	mem(45) := To_stdlogicvector(X"00");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"00");
	mem(49) := To_stdlogicvector(X"00");
	mem(50) := To_stdlogicvector(X"DD");
	mem(51) := To_stdlogicvector(X"BA");
	mem(52) := To_stdlogicvector(X"0D");
	mem(53) := To_stdlogicvector(X"60");
	mem(54) := To_stdlogicvector(X"AD");
	mem(55) := To_stdlogicvector(X"BB");
	mem(56) := To_stdlogicvector(X"AD");
	mem(57) := To_stdlogicvector(X"BB");
	mem(58) := To_stdlogicvector(X"DD");
	mem(59) := To_stdlogicvector(X"BA");
	mem(60) := To_stdlogicvector(X"AD");
	mem(61) := To_stdlogicvector(X"BB");
	mem(62) := To_stdlogicvector(X"AD");
	mem(63) := To_stdlogicvector(X"BB");
	mem(64) := To_stdlogicvector(X"AD");
	mem(65) := To_stdlogicvector(X"BB");
	mem(66) := To_stdlogicvector(X"AD");
	mem(67) := To_stdlogicvector(X"BB");
	mem(68) := To_stdlogicvector(X"AD");
	mem(69) := To_stdlogicvector(X"BB");
	mem(70) := To_stdlogicvector(X"AD");
	mem(71) := To_stdlogicvector(X"BB");
	mem(72) := To_stdlogicvector(X"AD");
	mem(73) := To_stdlogicvector(X"BB");
	mem(74) := To_stdlogicvector(X"AD");
	mem(75) := To_stdlogicvector(X"BB");
	mem(76) := To_stdlogicvector(X"AD");
	mem(77) := To_stdlogicvector(X"BB");
	mem(78) := To_stdlogicvector(X"AD");
	mem(79) := To_stdlogicvector(X"BB");
	mem(80) := To_stdlogicvector(X"AD");
	mem(81) := To_stdlogicvector(X"BB");
	mem(82) := To_stdlogicvector(X"AD");
	mem(83) := To_stdlogicvector(X"BB");
	mem(84) := To_stdlogicvector(X"AD");
	mem(85) := To_stdlogicvector(X"BB");
	mem(86) := To_stdlogicvector(X"AD");
	mem(87) := To_stdlogicvector(X"BB");
	mem(88) := To_stdlogicvector(X"AD");
	mem(89) := To_stdlogicvector(X"BB");
	mem(90) := To_stdlogicvector(X"AD");
	mem(91) := To_stdlogicvector(X"BB");
	mem(92) := To_stdlogicvector(X"AD");
	mem(93) := To_stdlogicvector(X"BB");
