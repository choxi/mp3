	mem(0) := To_stdlogicvector(X"03");
	mem(1) := To_stdlogicvector(X"E2");
	mem(2) := To_stdlogicvector(X"40");
	mem(3) := To_stdlogicvector(X"40");
	mem(4) := To_stdlogicvector(X"0F");
	mem(5) := To_stdlogicvector(X"6C");
	mem(6) := To_stdlogicvector(X"FE");
	mem(7) := To_stdlogicvector(X"0F");
	mem(8) := To_stdlogicvector(X"0C");
	mem(9) := To_stdlogicvector(X"6C");
	mem(10) := To_stdlogicvector(X"FE");
	mem(11) := To_stdlogicvector(X"0F");
	mem(12) := To_stdlogicvector(X"04");
	mem(13) := To_stdlogicvector(X"19");
	mem(14) := To_stdlogicvector(X"04");
	mem(15) := To_stdlogicvector(X"19");
	mem(16) := To_stdlogicvector(X"04");
	mem(17) := To_stdlogicvector(X"19");
	mem(18) := To_stdlogicvector(X"04");
	mem(19) := To_stdlogicvector(X"19");
	mem(20) := To_stdlogicvector(X"D0");
	mem(21) := To_stdlogicvector(X"BA");
	mem(22) := To_stdlogicvector(X"D1");
	mem(23) := To_stdlogicvector(X"BA");
	mem(24) := To_stdlogicvector(X"0D");
	mem(25) := To_stdlogicvector(X"60");
	mem(26) := To_stdlogicvector(X"D2");
	mem(27) := To_stdlogicvector(X"BA");
	mem(28) := To_stdlogicvector(X"D3");
	mem(29) := To_stdlogicvector(X"BA");
	mem(30) := To_stdlogicvector(X"DD");
	mem(31) := To_stdlogicvector(X"BA");
