	mem(0) := To_stdlogicvector(X"12");
	mem(1) := To_stdlogicvector(X"62");
	mem(2) := To_stdlogicvector(X"13");
	mem(3) := To_stdlogicvector(X"64");
	mem(4) := To_stdlogicvector(X"14");
	mem(5) := To_stdlogicvector(X"68");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"00");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"0D");
	mem(21) := To_stdlogicvector(X"0E");
	mem(22) := To_stdlogicvector(X"00");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"00");
	mem(25) := To_stdlogicvector(X"00");
	mem(26) := To_stdlogicvector(X"00");
	mem(27) := To_stdlogicvector(X"00");
	mem(28) := To_stdlogicvector(X"00");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"00");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"00");
	mem(33) := To_stdlogicvector(X"00");
	mem(34) := To_stdlogicvector(X"00");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"01");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"02");
	mem(39) := To_stdlogicvector(X"00");
	mem(40) := To_stdlogicvector(X"FF");
	mem(41) := To_stdlogicvector(X"FF");
	mem(42) := To_stdlogicvector(X"01");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"0D");
	mem(45) := To_stdlogicvector(X"60");
	mem(46) := To_stdlogicvector(X"DD");
	mem(47) := To_stdlogicvector(X"BA");
	mem(48) := To_stdlogicvector(X"42");
	mem(49) := To_stdlogicvector(X"16");
	mem(50) := To_stdlogicvector(X"82");
	mem(51) := To_stdlogicvector(X"5A");
	mem(52) := To_stdlogicvector(X"7F");
	mem(53) := To_stdlogicvector(X"9C");
	mem(54) := To_stdlogicvector(X"00");
	mem(55) := To_stdlogicvector(X"00");
	mem(56) := To_stdlogicvector(X"00");
	mem(57) := To_stdlogicvector(X"00");
	mem(58) := To_stdlogicvector(X"00");
	mem(59) := To_stdlogicvector(X"00");
	mem(60) := To_stdlogicvector(X"00");
	mem(61) := To_stdlogicvector(X"00");
	mem(62) := To_stdlogicvector(X"00");
	mem(63) := To_stdlogicvector(X"00");
	mem(64) := To_stdlogicvector(X"00");
	mem(65) := To_stdlogicvector(X"00");
	mem(66) := To_stdlogicvector(X"00");
	mem(67) := To_stdlogicvector(X"00");
	mem(68) := To_stdlogicvector(X"15");
	mem(69) := To_stdlogicvector(X"7C");
	mem(70) := To_stdlogicvector(X"15");
	mem(71) := To_stdlogicvector(X"6E");
	mem(72) := To_stdlogicvector(X"44");
	mem(73) := To_stdlogicvector(X"12");
	mem(74) := To_stdlogicvector(X"00");
	mem(75) := To_stdlogicvector(X"00");
	mem(76) := To_stdlogicvector(X"00");
	mem(77) := To_stdlogicvector(X"00");
	mem(78) := To_stdlogicvector(X"00");
	mem(79) := To_stdlogicvector(X"00");
	mem(80) := To_stdlogicvector(X"00");
	mem(81) := To_stdlogicvector(X"00");
	mem(82) := To_stdlogicvector(X"00");
	mem(83) := To_stdlogicvector(X"00");
	mem(84) := To_stdlogicvector(X"00");
	mem(85) := To_stdlogicvector(X"00");
	mem(86) := To_stdlogicvector(X"00");
	mem(87) := To_stdlogicvector(X"00");
	mem(88) := To_stdlogicvector(X"18");
	mem(89) := To_stdlogicvector(X"08");
	mem(90) := To_stdlogicvector(X"00");
	mem(91) := To_stdlogicvector(X"00");
	mem(92) := To_stdlogicvector(X"00");
	mem(93) := To_stdlogicvector(X"00");
	mem(94) := To_stdlogicvector(X"00");
	mem(95) := To_stdlogicvector(X"00");
	mem(96) := To_stdlogicvector(X"00");
	mem(97) := To_stdlogicvector(X"00");
	mem(98) := To_stdlogicvector(X"00");
	mem(99) := To_stdlogicvector(X"00");
	mem(100) := To_stdlogicvector(X"00");
	mem(101) := To_stdlogicvector(X"00");
	mem(102) := To_stdlogicvector(X"00");
	mem(103) := To_stdlogicvector(X"00");
	mem(104) := To_stdlogicvector(X"E3");
	mem(105) := To_stdlogicvector(X"0F");
	mem(106) := To_stdlogicvector(X"00");
	mem(107) := To_stdlogicvector(X"00");
	mem(108) := To_stdlogicvector(X"00");
	mem(109) := To_stdlogicvector(X"00");
	mem(110) := To_stdlogicvector(X"00");
	mem(111) := To_stdlogicvector(X"00");
	mem(112) := To_stdlogicvector(X"00");
	mem(113) := To_stdlogicvector(X"00");
	mem(114) := To_stdlogicvector(X"00");
	mem(115) := To_stdlogicvector(X"00");
	mem(116) := To_stdlogicvector(X"00");
	mem(117) := To_stdlogicvector(X"00");
	mem(118) := To_stdlogicvector(X"00");
	mem(119) := To_stdlogicvector(X"00");
	mem(120) := To_stdlogicvector(X"17");
	mem(121) := To_stdlogicvector(X"62");
	mem(122) := To_stdlogicvector(X"FE");
	mem(123) := To_stdlogicvector(X"0F");
	mem(124) := To_stdlogicvector(X"00");
	mem(125) := To_stdlogicvector(X"00");
	mem(126) := To_stdlogicvector(X"00");
	mem(127) := To_stdlogicvector(X"00");
	mem(128) := To_stdlogicvector(X"00");
	mem(129) := To_stdlogicvector(X"00");
	mem(130) := To_stdlogicvector(X"00");
	mem(131) := To_stdlogicvector(X"00");
	mem(132) := To_stdlogicvector(X"00");
	mem(133) := To_stdlogicvector(X"00");
	mem(134) := To_stdlogicvector(X"00");
	mem(135) := To_stdlogicvector(X"00");
	mem(136) := To_stdlogicvector(X"00");
	mem(137) := To_stdlogicvector(X"00");
	mem(138) := To_stdlogicvector(X"16");
	mem(139) := To_stdlogicvector(X"62");
	mem(140) := To_stdlogicvector(X"FE");
	mem(141) := To_stdlogicvector(X"0F");
	mem(142) := To_stdlogicvector(X"00");
	mem(143) := To_stdlogicvector(X"00");
	mem(144) := To_stdlogicvector(X"00");
	mem(145) := To_stdlogicvector(X"00");
	mem(146) := To_stdlogicvector(X"00");
	mem(147) := To_stdlogicvector(X"00");
	mem(148) := To_stdlogicvector(X"00");
	mem(149) := To_stdlogicvector(X"00");
	mem(150) := To_stdlogicvector(X"00");
	mem(151) := To_stdlogicvector(X"00");
	mem(152) := To_stdlogicvector(X"00");
	mem(153) := To_stdlogicvector(X"00");
	mem(154) := To_stdlogicvector(X"00");
	mem(155) := To_stdlogicvector(X"00");
