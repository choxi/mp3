	mem(0) := To_stdlogicvector(X"2F");
	mem(1) := To_stdlogicvector(X"12");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"0A");
	mem(13) := To_stdlogicvector(X"0E");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"00");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"D1");
	mem(25) := To_stdlogicvector(X"BA");
	mem(26) := To_stdlogicvector(X"D2");
	mem(27) := To_stdlogicvector(X"BA");
	mem(28) := To_stdlogicvector(X"D3");
	mem(29) := To_stdlogicvector(X"BA");
	mem(30) := To_stdlogicvector(X"D4");
	mem(31) := To_stdlogicvector(X"BA");
	mem(32) := To_stdlogicvector(X"D5");
	mem(33) := To_stdlogicvector(X"BA");
	mem(34) := To_stdlogicvector(X"3F");
	mem(35) := To_stdlogicvector(X"12");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"00");
	mem(39) := To_stdlogicvector(X"00");
	mem(40) := To_stdlogicvector(X"00");
	mem(41) := To_stdlogicvector(X"00");
	mem(42) := To_stdlogicvector(X"00");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"00");
	mem(45) := To_stdlogicvector(X"00");
	mem(46) := To_stdlogicvector(X"0A");
	mem(47) := To_stdlogicvector(X"08");
	mem(48) := To_stdlogicvector(X"00");
	mem(49) := To_stdlogicvector(X"00");
	mem(50) := To_stdlogicvector(X"00");
	mem(51) := To_stdlogicvector(X"00");
	mem(52) := To_stdlogicvector(X"00");
	mem(53) := To_stdlogicvector(X"00");
	mem(54) := To_stdlogicvector(X"00");
	mem(55) := To_stdlogicvector(X"00");
	mem(56) := To_stdlogicvector(X"00");
	mem(57) := To_stdlogicvector(X"00");
	mem(58) := To_stdlogicvector(X"D1");
	mem(59) := To_stdlogicvector(X"BA");
	mem(60) := To_stdlogicvector(X"D2");
	mem(61) := To_stdlogicvector(X"BA");
	mem(62) := To_stdlogicvector(X"D3");
	mem(63) := To_stdlogicvector(X"BA");
	mem(64) := To_stdlogicvector(X"D4");
	mem(65) := To_stdlogicvector(X"BA");
	mem(66) := To_stdlogicvector(X"D5");
	mem(67) := To_stdlogicvector(X"BA");
	mem(68) := To_stdlogicvector(X"20");
	mem(69) := To_stdlogicvector(X"12");
	mem(70) := To_stdlogicvector(X"00");
	mem(71) := To_stdlogicvector(X"00");
	mem(72) := To_stdlogicvector(X"00");
	mem(73) := To_stdlogicvector(X"00");
	mem(74) := To_stdlogicvector(X"00");
	mem(75) := To_stdlogicvector(X"00");
	mem(76) := To_stdlogicvector(X"00");
	mem(77) := To_stdlogicvector(X"00");
	mem(78) := To_stdlogicvector(X"00");
	mem(79) := To_stdlogicvector(X"00");
	mem(80) := To_stdlogicvector(X"0A");
	mem(81) := To_stdlogicvector(X"04");
	mem(82) := To_stdlogicvector(X"00");
	mem(83) := To_stdlogicvector(X"00");
	mem(84) := To_stdlogicvector(X"00");
	mem(85) := To_stdlogicvector(X"00");
	mem(86) := To_stdlogicvector(X"00");
	mem(87) := To_stdlogicvector(X"00");
	mem(88) := To_stdlogicvector(X"00");
	mem(89) := To_stdlogicvector(X"00");
	mem(90) := To_stdlogicvector(X"00");
	mem(91) := To_stdlogicvector(X"00");
	mem(92) := To_stdlogicvector(X"D1");
	mem(93) := To_stdlogicvector(X"BA");
	mem(94) := To_stdlogicvector(X"D2");
	mem(95) := To_stdlogicvector(X"BA");
	mem(96) := To_stdlogicvector(X"D3");
	mem(97) := To_stdlogicvector(X"BA");
	mem(98) := To_stdlogicvector(X"D4");
	mem(99) := To_stdlogicvector(X"BA");
	mem(100) := To_stdlogicvector(X"D5");
	mem(101) := To_stdlogicvector(X"BA");
	mem(102) := To_stdlogicvector(X"27");
	mem(103) := To_stdlogicvector(X"12");
	mem(104) := To_stdlogicvector(X"00");
	mem(105) := To_stdlogicvector(X"00");
	mem(106) := To_stdlogicvector(X"00");
	mem(107) := To_stdlogicvector(X"00");
	mem(108) := To_stdlogicvector(X"00");
	mem(109) := To_stdlogicvector(X"00");
	mem(110) := To_stdlogicvector(X"00");
	mem(111) := To_stdlogicvector(X"00");
	mem(112) := To_stdlogicvector(X"00");
	mem(113) := To_stdlogicvector(X"00");
	mem(114) := To_stdlogicvector(X"0A");
	mem(115) := To_stdlogicvector(X"02");
	mem(116) := To_stdlogicvector(X"00");
	mem(117) := To_stdlogicvector(X"00");
	mem(118) := To_stdlogicvector(X"00");
	mem(119) := To_stdlogicvector(X"00");
	mem(120) := To_stdlogicvector(X"00");
	mem(121) := To_stdlogicvector(X"00");
	mem(122) := To_stdlogicvector(X"00");
	mem(123) := To_stdlogicvector(X"00");
	mem(124) := To_stdlogicvector(X"00");
	mem(125) := To_stdlogicvector(X"00");
	mem(126) := To_stdlogicvector(X"D1");
	mem(127) := To_stdlogicvector(X"BA");
	mem(128) := To_stdlogicvector(X"D2");
	mem(129) := To_stdlogicvector(X"BA");
	mem(130) := To_stdlogicvector(X"D3");
	mem(131) := To_stdlogicvector(X"BA");
	mem(132) := To_stdlogicvector(X"D4");
	mem(133) := To_stdlogicvector(X"BA");
	mem(134) := To_stdlogicvector(X"D5");
	mem(135) := To_stdlogicvector(X"BA");
	mem(136) := To_stdlogicvector(X"3F");
	mem(137) := To_stdlogicvector(X"12");
	mem(138) := To_stdlogicvector(X"00");
	mem(139) := To_stdlogicvector(X"00");
	mem(140) := To_stdlogicvector(X"00");
	mem(141) := To_stdlogicvector(X"00");
	mem(142) := To_stdlogicvector(X"00");
	mem(143) := To_stdlogicvector(X"00");
	mem(144) := To_stdlogicvector(X"00");
	mem(145) := To_stdlogicvector(X"00");
	mem(146) := To_stdlogicvector(X"00");
	mem(147) := To_stdlogicvector(X"00");
	mem(148) := To_stdlogicvector(X"0A");
	mem(149) := To_stdlogicvector(X"0C");
	mem(150) := To_stdlogicvector(X"00");
	mem(151) := To_stdlogicvector(X"00");
	mem(152) := To_stdlogicvector(X"00");
	mem(153) := To_stdlogicvector(X"00");
	mem(154) := To_stdlogicvector(X"00");
	mem(155) := To_stdlogicvector(X"00");
	mem(156) := To_stdlogicvector(X"00");
	mem(157) := To_stdlogicvector(X"00");
	mem(158) := To_stdlogicvector(X"00");
	mem(159) := To_stdlogicvector(X"00");
	mem(160) := To_stdlogicvector(X"D1");
	mem(161) := To_stdlogicvector(X"BA");
	mem(162) := To_stdlogicvector(X"D2");
	mem(163) := To_stdlogicvector(X"BA");
	mem(164) := To_stdlogicvector(X"D3");
	mem(165) := To_stdlogicvector(X"BA");
	mem(166) := To_stdlogicvector(X"D4");
	mem(167) := To_stdlogicvector(X"BA");
	mem(168) := To_stdlogicvector(X"D5");
	mem(169) := To_stdlogicvector(X"BA");
	mem(170) := To_stdlogicvector(X"20");
	mem(171) := To_stdlogicvector(X"12");
	mem(172) := To_stdlogicvector(X"00");
	mem(173) := To_stdlogicvector(X"00");
	mem(174) := To_stdlogicvector(X"00");
	mem(175) := To_stdlogicvector(X"00");
	mem(176) := To_stdlogicvector(X"00");
	mem(177) := To_stdlogicvector(X"00");
	mem(178) := To_stdlogicvector(X"00");
	mem(179) := To_stdlogicvector(X"00");
	mem(180) := To_stdlogicvector(X"00");
	mem(181) := To_stdlogicvector(X"00");
	mem(182) := To_stdlogicvector(X"0A");
	mem(183) := To_stdlogicvector(X"0C");
	mem(184) := To_stdlogicvector(X"00");
	mem(185) := To_stdlogicvector(X"00");
	mem(186) := To_stdlogicvector(X"00");
	mem(187) := To_stdlogicvector(X"00");
	mem(188) := To_stdlogicvector(X"00");
	mem(189) := To_stdlogicvector(X"00");
	mem(190) := To_stdlogicvector(X"00");
	mem(191) := To_stdlogicvector(X"00");
	mem(192) := To_stdlogicvector(X"00");
	mem(193) := To_stdlogicvector(X"00");
	mem(194) := To_stdlogicvector(X"D1");
	mem(195) := To_stdlogicvector(X"BA");
	mem(196) := To_stdlogicvector(X"D2");
	mem(197) := To_stdlogicvector(X"BA");
	mem(198) := To_stdlogicvector(X"D3");
	mem(199) := To_stdlogicvector(X"BA");
	mem(200) := To_stdlogicvector(X"D4");
	mem(201) := To_stdlogicvector(X"BA");
	mem(202) := To_stdlogicvector(X"D5");
	mem(203) := To_stdlogicvector(X"BA");
	mem(204) := To_stdlogicvector(X"32");
	mem(205) := To_stdlogicvector(X"12");
	mem(206) := To_stdlogicvector(X"00");
	mem(207) := To_stdlogicvector(X"00");
	mem(208) := To_stdlogicvector(X"00");
	mem(209) := To_stdlogicvector(X"00");
	mem(210) := To_stdlogicvector(X"00");
	mem(211) := To_stdlogicvector(X"00");
	mem(212) := To_stdlogicvector(X"00");
	mem(213) := To_stdlogicvector(X"00");
	mem(214) := To_stdlogicvector(X"00");
	mem(215) := To_stdlogicvector(X"00");
	mem(216) := To_stdlogicvector(X"0A");
	mem(217) := To_stdlogicvector(X"0A");
	mem(218) := To_stdlogicvector(X"00");
	mem(219) := To_stdlogicvector(X"00");
	mem(220) := To_stdlogicvector(X"00");
	mem(221) := To_stdlogicvector(X"00");
	mem(222) := To_stdlogicvector(X"00");
	mem(223) := To_stdlogicvector(X"00");
	mem(224) := To_stdlogicvector(X"00");
	mem(225) := To_stdlogicvector(X"00");
	mem(226) := To_stdlogicvector(X"00");
	mem(227) := To_stdlogicvector(X"00");
	mem(228) := To_stdlogicvector(X"D1");
	mem(229) := To_stdlogicvector(X"BA");
	mem(230) := To_stdlogicvector(X"D2");
	mem(231) := To_stdlogicvector(X"BA");
	mem(232) := To_stdlogicvector(X"D3");
	mem(233) := To_stdlogicvector(X"BA");
	mem(234) := To_stdlogicvector(X"D4");
	mem(235) := To_stdlogicvector(X"BA");
	mem(236) := To_stdlogicvector(X"D5");
	mem(237) := To_stdlogicvector(X"BA");
	mem(238) := To_stdlogicvector(X"29");
	mem(239) := To_stdlogicvector(X"12");
	mem(240) := To_stdlogicvector(X"00");
	mem(241) := To_stdlogicvector(X"00");
	mem(242) := To_stdlogicvector(X"00");
	mem(243) := To_stdlogicvector(X"00");
	mem(244) := To_stdlogicvector(X"00");
	mem(245) := To_stdlogicvector(X"00");
	mem(246) := To_stdlogicvector(X"00");
	mem(247) := To_stdlogicvector(X"00");
	mem(248) := To_stdlogicvector(X"00");
	mem(249) := To_stdlogicvector(X"00");
	mem(250) := To_stdlogicvector(X"0A");
	mem(251) := To_stdlogicvector(X"0A");
	mem(252) := To_stdlogicvector(X"00");
	mem(253) := To_stdlogicvector(X"00");
	mem(254) := To_stdlogicvector(X"00");
	mem(255) := To_stdlogicvector(X"00");
	mem(256) := To_stdlogicvector(X"00");
	mem(257) := To_stdlogicvector(X"00");
	mem(258) := To_stdlogicvector(X"00");
	mem(259) := To_stdlogicvector(X"00");
	mem(260) := To_stdlogicvector(X"00");
	mem(261) := To_stdlogicvector(X"00");
	mem(262) := To_stdlogicvector(X"D1");
	mem(263) := To_stdlogicvector(X"BA");
	mem(264) := To_stdlogicvector(X"D2");
	mem(265) := To_stdlogicvector(X"BA");
	mem(266) := To_stdlogicvector(X"D3");
	mem(267) := To_stdlogicvector(X"BA");
	mem(268) := To_stdlogicvector(X"D4");
	mem(269) := To_stdlogicvector(X"BA");
	mem(270) := To_stdlogicvector(X"D5");
	mem(271) := To_stdlogicvector(X"BA");
	mem(272) := To_stdlogicvector(X"20");
	mem(273) := To_stdlogicvector(X"12");
	mem(274) := To_stdlogicvector(X"00");
	mem(275) := To_stdlogicvector(X"00");
	mem(276) := To_stdlogicvector(X"00");
	mem(277) := To_stdlogicvector(X"00");
	mem(278) := To_stdlogicvector(X"00");
	mem(279) := To_stdlogicvector(X"00");
	mem(280) := To_stdlogicvector(X"00");
	mem(281) := To_stdlogicvector(X"00");
	mem(282) := To_stdlogicvector(X"00");
	mem(283) := To_stdlogicvector(X"00");
	mem(284) := To_stdlogicvector(X"0A");
	mem(285) := To_stdlogicvector(X"06");
	mem(286) := To_stdlogicvector(X"00");
	mem(287) := To_stdlogicvector(X"00");
	mem(288) := To_stdlogicvector(X"00");
	mem(289) := To_stdlogicvector(X"00");
	mem(290) := To_stdlogicvector(X"00");
	mem(291) := To_stdlogicvector(X"00");
	mem(292) := To_stdlogicvector(X"00");
	mem(293) := To_stdlogicvector(X"00");
	mem(294) := To_stdlogicvector(X"00");
	mem(295) := To_stdlogicvector(X"00");
	mem(296) := To_stdlogicvector(X"D1");
	mem(297) := To_stdlogicvector(X"BA");
	mem(298) := To_stdlogicvector(X"D2");
	mem(299) := To_stdlogicvector(X"BA");
	mem(300) := To_stdlogicvector(X"D3");
	mem(301) := To_stdlogicvector(X"BA");
	mem(302) := To_stdlogicvector(X"D4");
	mem(303) := To_stdlogicvector(X"BA");
	mem(304) := To_stdlogicvector(X"D5");
	mem(305) := To_stdlogicvector(X"BA");
	mem(306) := To_stdlogicvector(X"2B");
	mem(307) := To_stdlogicvector(X"12");
	mem(308) := To_stdlogicvector(X"00");
	mem(309) := To_stdlogicvector(X"00");
	mem(310) := To_stdlogicvector(X"00");
	mem(311) := To_stdlogicvector(X"00");
	mem(312) := To_stdlogicvector(X"00");
	mem(313) := To_stdlogicvector(X"00");
	mem(314) := To_stdlogicvector(X"00");
	mem(315) := To_stdlogicvector(X"00");
	mem(316) := To_stdlogicvector(X"00");
	mem(317) := To_stdlogicvector(X"00");
	mem(318) := To_stdlogicvector(X"0A");
	mem(319) := To_stdlogicvector(X"06");
	mem(320) := To_stdlogicvector(X"00");
	mem(321) := To_stdlogicvector(X"00");
	mem(322) := To_stdlogicvector(X"00");
	mem(323) := To_stdlogicvector(X"00");
	mem(324) := To_stdlogicvector(X"00");
	mem(325) := To_stdlogicvector(X"00");
	mem(326) := To_stdlogicvector(X"00");
	mem(327) := To_stdlogicvector(X"00");
	mem(328) := To_stdlogicvector(X"00");
	mem(329) := To_stdlogicvector(X"00");
	mem(330) := To_stdlogicvector(X"D1");
	mem(331) := To_stdlogicvector(X"BA");
	mem(332) := To_stdlogicvector(X"D2");
	mem(333) := To_stdlogicvector(X"BA");
	mem(334) := To_stdlogicvector(X"D3");
	mem(335) := To_stdlogicvector(X"BA");
	mem(336) := To_stdlogicvector(X"D4");
	mem(337) := To_stdlogicvector(X"BA");
	mem(338) := To_stdlogicvector(X"D5");
	mem(339) := To_stdlogicvector(X"BA");
	mem(340) := To_stdlogicvector(X"00");
	mem(341) := To_stdlogicvector(X"00");
	mem(342) := To_stdlogicvector(X"00");
	mem(343) := To_stdlogicvector(X"00");
	mem(344) := To_stdlogicvector(X"00");
	mem(345) := To_stdlogicvector(X"00");
	mem(346) := To_stdlogicvector(X"00");
	mem(347) := To_stdlogicvector(X"00");
	mem(348) := To_stdlogicvector(X"00");
	mem(349) := To_stdlogicvector(X"00");
	mem(350) := To_stdlogicvector(X"FA");
	mem(351) := To_stdlogicvector(X"0F");
	mem(352) := To_stdlogicvector(X"00");
	mem(353) := To_stdlogicvector(X"00");
	mem(354) := To_stdlogicvector(X"00");
	mem(355) := To_stdlogicvector(X"00");
	mem(356) := To_stdlogicvector(X"00");
	mem(357) := To_stdlogicvector(X"00");
	mem(358) := To_stdlogicvector(X"00");
	mem(359) := To_stdlogicvector(X"00");
	mem(360) := To_stdlogicvector(X"00");
	mem(361) := To_stdlogicvector(X"00");
	mem(362) := To_stdlogicvector(X"DD");
	mem(363) := To_stdlogicvector(X"BA");
