	mem(0) := To_stdlogicvector(X"61");
	mem(1) := To_stdlogicvector(X"12");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"FA");
	mem(13) := To_stdlogicvector(X"0F");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
