	mem(40) := To_stdlogicvector(X"1E");
	mem(41) := To_stdlogicvector(X"F0");
	mem(42) := To_stdlogicvector(X"13");
	mem(43) := To_stdlogicvector(X"E2");
	mem(44) := To_stdlogicvector(X"40");
	mem(45) := To_stdlogicvector(X"C0");
	mem(46) := To_stdlogicvector(X"21");
	mem(47) := To_stdlogicvector(X"10");
	mem(48) := To_stdlogicvector(X"21");
	mem(49) := To_stdlogicvector(X"10");
	mem(50) := To_stdlogicvector(X"21");
	mem(51) := To_stdlogicvector(X"10");
	mem(52) := To_stdlogicvector(X"21");
	mem(53) := To_stdlogicvector(X"10");
	mem(54) := To_stdlogicvector(X"21");
	mem(55) := To_stdlogicvector(X"10");
	mem(56) := To_stdlogicvector(X"21");
	mem(57) := To_stdlogicvector(X"10");
	mem(58) := To_stdlogicvector(X"21");
	mem(59) := To_stdlogicvector(X"10");
	mem(60) := To_stdlogicvector(X"4E");
	mem(61) := To_stdlogicvector(X"00");
	mem(62) := To_stdlogicvector(X"21");
	mem(63) := To_stdlogicvector(X"10");
	mem(64) := To_stdlogicvector(X"21");
	mem(65) := To_stdlogicvector(X"10");
	mem(66) := To_stdlogicvector(X"21");
	mem(67) := To_stdlogicvector(X"10");
	mem(68) := To_stdlogicvector(X"21");
	mem(69) := To_stdlogicvector(X"10");
	mem(70) := To_stdlogicvector(X"21");
	mem(71) := To_stdlogicvector(X"10");
	mem(72) := To_stdlogicvector(X"21");
	mem(73) := To_stdlogicvector(X"10");
	mem(74) := To_stdlogicvector(X"21");
	mem(75) := To_stdlogicvector(X"10");
	mem(76) := To_stdlogicvector(X"21");
	mem(77) := To_stdlogicvector(X"10");
	mem(78) := To_stdlogicvector(X"2F");
	mem(79) := To_stdlogicvector(X"19");
	mem(80) := To_stdlogicvector(X"C0");
	mem(81) := To_stdlogicvector(X"C1");
	mem(82) := To_stdlogicvector(X"FF");
	mem(83) := To_stdlogicvector(X"0F");
