	mem(0) := To_stdlogicvector(X"07");
	mem(1) := To_stdlogicvector(X"0E");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"00");
	mem(14) := To_stdlogicvector(X"80");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"07");
	mem(17) := To_stdlogicvector(X"60");
	mem(18) := To_stdlogicvector(X"00");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"00");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"00");
	mem(25) := To_stdlogicvector(X"00");
	mem(26) := To_stdlogicvector(X"00");
	mem(27) := To_stdlogicvector(X"00");
	mem(28) := To_stdlogicvector(X"06");
	mem(29) := To_stdlogicvector(X"62");
	mem(30) := To_stdlogicvector(X"08");
	mem(31) := To_stdlogicvector(X"66");
	mem(32) := To_stdlogicvector(X"07");
	mem(33) := To_stdlogicvector(X"64");
	mem(34) := To_stdlogicvector(X"09");
	mem(35) := To_stdlogicvector(X"68");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"09");
	mem(39) := To_stdlogicvector(X"72");
	mem(40) := To_stdlogicvector(X"08");
	mem(41) := To_stdlogicvector(X"74");
	mem(42) := To_stdlogicvector(X"07");
	mem(43) := To_stdlogicvector(X"76");
	mem(44) := To_stdlogicvector(X"06");
	mem(45) := To_stdlogicvector(X"78");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"06");
	mem(49) := To_stdlogicvector(X"62");
	mem(50) := To_stdlogicvector(X"07");
	mem(51) := To_stdlogicvector(X"64");
	mem(52) := To_stdlogicvector(X"08");
	mem(53) := To_stdlogicvector(X"66");
	mem(54) := To_stdlogicvector(X"09");
	mem(55) := To_stdlogicvector(X"68");
	mem(56) := To_stdlogicvector(X"12");
	mem(57) := To_stdlogicvector(X"0E");
	mem(58) := To_stdlogicvector(X"00");
	mem(59) := To_stdlogicvector(X"00");
	mem(60) := To_stdlogicvector(X"00");
	mem(61) := To_stdlogicvector(X"00");
	mem(62) := To_stdlogicvector(X"00");
	mem(63) := To_stdlogicvector(X"00");
	mem(64) := To_stdlogicvector(X"00");
	mem(65) := To_stdlogicvector(X"00");
	mem(66) := To_stdlogicvector(X"00");
	mem(67) := To_stdlogicvector(X"00");
	mem(68) := To_stdlogicvector(X"00");
	mem(69) := To_stdlogicvector(X"00");
	mem(70) := To_stdlogicvector(X"00");
	mem(71) := To_stdlogicvector(X"00");
	mem(72) := To_stdlogicvector(X"00");
	mem(73) := To_stdlogicvector(X"00");
	mem(74) := To_stdlogicvector(X"00");
	mem(75) := To_stdlogicvector(X"00");
	mem(76) := To_stdlogicvector(X"00");
	mem(77) := To_stdlogicvector(X"00");
	mem(78) := To_stdlogicvector(X"00");
	mem(79) := To_stdlogicvector(X"00");
	mem(80) := To_stdlogicvector(X"00");
	mem(81) := To_stdlogicvector(X"00");
	mem(82) := To_stdlogicvector(X"00");
	mem(83) := To_stdlogicvector(X"00");
	mem(84) := To_stdlogicvector(X"00");
	mem(85) := To_stdlogicvector(X"00");
	mem(86) := To_stdlogicvector(X"00");
	mem(87) := To_stdlogicvector(X"00");
	mem(88) := To_stdlogicvector(X"00");
	mem(89) := To_stdlogicvector(X"00");
	mem(90) := To_stdlogicvector(X"00");
	mem(91) := To_stdlogicvector(X"00");
	mem(92) := To_stdlogicvector(X"00");
	mem(93) := To_stdlogicvector(X"00");
	mem(94) := To_stdlogicvector(X"42");
	mem(95) := To_stdlogicvector(X"1A");
	mem(96) := To_stdlogicvector(X"C4");
	mem(97) := To_stdlogicvector(X"1C");
	mem(98) := To_stdlogicvector(X"00");
	mem(99) := To_stdlogicvector(X"00");
	mem(100) := To_stdlogicvector(X"00");
	mem(101) := To_stdlogicvector(X"00");
	mem(102) := To_stdlogicvector(X"00");
	mem(103) := To_stdlogicvector(X"00");
	mem(104) := To_stdlogicvector(X"00");
	mem(105) := To_stdlogicvector(X"00");
	mem(106) := To_stdlogicvector(X"18");
	mem(107) := To_stdlogicvector(X"7A");
	mem(108) := To_stdlogicvector(X"46");
	mem(109) := To_stdlogicvector(X"1F");
	mem(110) := To_stdlogicvector(X"00");
	mem(111) := To_stdlogicvector(X"00");
	mem(112) := To_stdlogicvector(X"00");
	mem(113) := To_stdlogicvector(X"00");
	mem(114) := To_stdlogicvector(X"00");
	mem(115) := To_stdlogicvector(X"00");
	mem(116) := To_stdlogicvector(X"00");
	mem(117) := To_stdlogicvector(X"00");
	mem(118) := To_stdlogicvector(X"10");
	mem(119) := To_stdlogicvector(X"7E");
	mem(120) := To_stdlogicvector(X"10");
	mem(121) := To_stdlogicvector(X"62");
	mem(122) := To_stdlogicvector(X"FF");
	mem(123) := To_stdlogicvector(X"0F");
	mem(124) := To_stdlogicvector(X"00");
	mem(125) := To_stdlogicvector(X"00");
	mem(126) := To_stdlogicvector(X"00");
	mem(127) := To_stdlogicvector(X"00");
	mem(128) := To_stdlogicvector(X"00");
	mem(129) := To_stdlogicvector(X"00");
	mem(130) := To_stdlogicvector(X"00");
	mem(131) := To_stdlogicvector(X"00");
	mem(132) := To_stdlogicvector(X"00");
	mem(133) := To_stdlogicvector(X"00");
	mem(134) := To_stdlogicvector(X"00");
	mem(135) := To_stdlogicvector(X"00");
	mem(136) := To_stdlogicvector(X"00");
	mem(137) := To_stdlogicvector(X"00");
	mem(138) := To_stdlogicvector(X"00");
	mem(139) := To_stdlogicvector(X"00");
	mem(140) := To_stdlogicvector(X"09");
	mem(141) := To_stdlogicvector(X"00");
	mem(142) := To_stdlogicvector(X"02");
	mem(143) := To_stdlogicvector(X"00");
	mem(144) := To_stdlogicvector(X"01");
	mem(145) := To_stdlogicvector(X"00");
	mem(146) := To_stdlogicvector(X"03");
	mem(147) := To_stdlogicvector(X"00");
	mem(148) := To_stdlogicvector(X"00");
	mem(149) := To_stdlogicvector(X"00");
	mem(150) := To_stdlogicvector(X"00");
	mem(151) := To_stdlogicvector(X"00");
	mem(152) := To_stdlogicvector(X"00");
	mem(153) := To_stdlogicvector(X"00");
	mem(154) := To_stdlogicvector(X"00");
	mem(155) := To_stdlogicvector(X"00");
	mem(156) := To_stdlogicvector(X"00");
	mem(157) := To_stdlogicvector(X"00");
	mem(158) := To_stdlogicvector(X"00");
	mem(159) := To_stdlogicvector(X"00");
	mem(160) := To_stdlogicvector(X"00");
	mem(161) := To_stdlogicvector(X"00");
	mem(162) := To_stdlogicvector(X"00");
	mem(163) := To_stdlogicvector(X"00");
	mem(164) := To_stdlogicvector(X"00");
	mem(165) := To_stdlogicvector(X"00");
	mem(166) := To_stdlogicvector(X"00");
	mem(167) := To_stdlogicvector(X"00");
	mem(168) := To_stdlogicvector(X"00");
	mem(169) := To_stdlogicvector(X"00");
	mem(170) := To_stdlogicvector(X"00");
	mem(171) := To_stdlogicvector(X"00");
	mem(172) := To_stdlogicvector(X"00");
	mem(173) := To_stdlogicvector(X"00");
	mem(174) := To_stdlogicvector(X"00");
	mem(175) := To_stdlogicvector(X"00");
	mem(176) := To_stdlogicvector(X"00");
	mem(177) := To_stdlogicvector(X"00");
	mem(178) := To_stdlogicvector(X"00");
	mem(179) := To_stdlogicvector(X"00");
	mem(180) := To_stdlogicvector(X"00");
	mem(181) := To_stdlogicvector(X"00");
	mem(182) := To_stdlogicvector(X"00");
	mem(183) := To_stdlogicvector(X"00");
	mem(184) := To_stdlogicvector(X"00");
	mem(185) := To_stdlogicvector(X"00");
	mem(186) := To_stdlogicvector(X"00");
	mem(187) := To_stdlogicvector(X"00");
	mem(188) := To_stdlogicvector(X"00");
	mem(189) := To_stdlogicvector(X"00");
	mem(190) := To_stdlogicvector(X"00");
	mem(191) := To_stdlogicvector(X"00");
