	mem(0) := To_stdlogicvector(X"2F");
	mem(1) := To_stdlogicvector(X"12");
	mem(2) := To_stdlogicvector(X"0B");
	mem(3) := To_stdlogicvector(X"08");
	mem(4) := To_stdlogicvector(X"67");
	mem(5) := To_stdlogicvector(X"14");
	mem(6) := To_stdlogicvector(X"28");
	mem(7) := To_stdlogicvector(X"16");
	mem(8) := To_stdlogicvector(X"29");
	mem(9) := To_stdlogicvector(X"18");
	mem(10) := To_stdlogicvector(X"2A");
	mem(11) := To_stdlogicvector(X"1A");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"00");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"D1");
	mem(17) := To_stdlogicvector(X"BA");
	mem(18) := To_stdlogicvector(X"D2");
	mem(19) := To_stdlogicvector(X"BA");
	mem(20) := To_stdlogicvector(X"D3");
	mem(21) := To_stdlogicvector(X"BA");
	mem(22) := To_stdlogicvector(X"D4");
	mem(23) := To_stdlogicvector(X"BA");
	mem(24) := To_stdlogicvector(X"D5");
	mem(25) := To_stdlogicvector(X"BA");
	mem(26) := To_stdlogicvector(X"3F");
	mem(27) := To_stdlogicvector(X"12");
	mem(28) := To_stdlogicvector(X"00");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"00");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"00");
	mem(33) := To_stdlogicvector(X"00");
	mem(34) := To_stdlogicvector(X"00");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"00");
	mem(37) := To_stdlogicvector(X"00");
	mem(38) := To_stdlogicvector(X"0A");
	mem(39) := To_stdlogicvector(X"08");
	mem(40) := To_stdlogicvector(X"00");
	mem(41) := To_stdlogicvector(X"00");
	mem(42) := To_stdlogicvector(X"00");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"00");
	mem(45) := To_stdlogicvector(X"00");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"00");
	mem(49) := To_stdlogicvector(X"00");
	mem(50) := To_stdlogicvector(X"D1");
	mem(51) := To_stdlogicvector(X"BA");
	mem(52) := To_stdlogicvector(X"D2");
	mem(53) := To_stdlogicvector(X"BA");
	mem(54) := To_stdlogicvector(X"D3");
	mem(55) := To_stdlogicvector(X"BA");
	mem(56) := To_stdlogicvector(X"D4");
	mem(57) := To_stdlogicvector(X"BA");
	mem(58) := To_stdlogicvector(X"D5");
	mem(59) := To_stdlogicvector(X"BA");
	mem(60) := To_stdlogicvector(X"20");
	mem(61) := To_stdlogicvector(X"12");
	mem(62) := To_stdlogicvector(X"00");
	mem(63) := To_stdlogicvector(X"00");
	mem(64) := To_stdlogicvector(X"00");
	mem(65) := To_stdlogicvector(X"00");
	mem(66) := To_stdlogicvector(X"00");
	mem(67) := To_stdlogicvector(X"00");
	mem(68) := To_stdlogicvector(X"00");
	mem(69) := To_stdlogicvector(X"00");
	mem(70) := To_stdlogicvector(X"00");
	mem(71) := To_stdlogicvector(X"00");
	mem(72) := To_stdlogicvector(X"0A");
	mem(73) := To_stdlogicvector(X"04");
	mem(74) := To_stdlogicvector(X"00");
	mem(75) := To_stdlogicvector(X"00");
	mem(76) := To_stdlogicvector(X"00");
	mem(77) := To_stdlogicvector(X"00");
	mem(78) := To_stdlogicvector(X"00");
	mem(79) := To_stdlogicvector(X"00");
	mem(80) := To_stdlogicvector(X"00");
	mem(81) := To_stdlogicvector(X"00");
	mem(82) := To_stdlogicvector(X"00");
	mem(83) := To_stdlogicvector(X"00");
	mem(84) := To_stdlogicvector(X"D1");
	mem(85) := To_stdlogicvector(X"BA");
	mem(86) := To_stdlogicvector(X"D2");
	mem(87) := To_stdlogicvector(X"BA");
	mem(88) := To_stdlogicvector(X"D3");
	mem(89) := To_stdlogicvector(X"BA");
	mem(90) := To_stdlogicvector(X"D4");
	mem(91) := To_stdlogicvector(X"BA");
	mem(92) := To_stdlogicvector(X"D5");
	mem(93) := To_stdlogicvector(X"BA");
	mem(94) := To_stdlogicvector(X"27");
	mem(95) := To_stdlogicvector(X"12");
	mem(96) := To_stdlogicvector(X"00");
	mem(97) := To_stdlogicvector(X"00");
	mem(98) := To_stdlogicvector(X"00");
	mem(99) := To_stdlogicvector(X"00");
	mem(100) := To_stdlogicvector(X"00");
	mem(101) := To_stdlogicvector(X"00");
	mem(102) := To_stdlogicvector(X"00");
	mem(103) := To_stdlogicvector(X"00");
	mem(104) := To_stdlogicvector(X"00");
	mem(105) := To_stdlogicvector(X"00");
	mem(106) := To_stdlogicvector(X"0A");
	mem(107) := To_stdlogicvector(X"02");
	mem(108) := To_stdlogicvector(X"00");
	mem(109) := To_stdlogicvector(X"00");
	mem(110) := To_stdlogicvector(X"00");
	mem(111) := To_stdlogicvector(X"00");
	mem(112) := To_stdlogicvector(X"00");
	mem(113) := To_stdlogicvector(X"00");
	mem(114) := To_stdlogicvector(X"00");
	mem(115) := To_stdlogicvector(X"00");
	mem(116) := To_stdlogicvector(X"00");
	mem(117) := To_stdlogicvector(X"00");
	mem(118) := To_stdlogicvector(X"D1");
	mem(119) := To_stdlogicvector(X"BA");
	mem(120) := To_stdlogicvector(X"D2");
	mem(121) := To_stdlogicvector(X"BA");
	mem(122) := To_stdlogicvector(X"D3");
	mem(123) := To_stdlogicvector(X"BA");
	mem(124) := To_stdlogicvector(X"D4");
	mem(125) := To_stdlogicvector(X"BA");
	mem(126) := To_stdlogicvector(X"D5");
	mem(127) := To_stdlogicvector(X"BA");
	mem(128) := To_stdlogicvector(X"3F");
	mem(129) := To_stdlogicvector(X"12");
	mem(130) := To_stdlogicvector(X"00");
	mem(131) := To_stdlogicvector(X"00");
	mem(132) := To_stdlogicvector(X"00");
	mem(133) := To_stdlogicvector(X"00");
	mem(134) := To_stdlogicvector(X"00");
	mem(135) := To_stdlogicvector(X"00");
	mem(136) := To_stdlogicvector(X"00");
	mem(137) := To_stdlogicvector(X"00");
	mem(138) := To_stdlogicvector(X"00");
	mem(139) := To_stdlogicvector(X"00");
	mem(140) := To_stdlogicvector(X"0A");
	mem(141) := To_stdlogicvector(X"0C");
	mem(142) := To_stdlogicvector(X"00");
	mem(143) := To_stdlogicvector(X"00");
	mem(144) := To_stdlogicvector(X"00");
	mem(145) := To_stdlogicvector(X"00");
	mem(146) := To_stdlogicvector(X"00");
	mem(147) := To_stdlogicvector(X"00");
	mem(148) := To_stdlogicvector(X"00");
	mem(149) := To_stdlogicvector(X"00");
	mem(150) := To_stdlogicvector(X"00");
	mem(151) := To_stdlogicvector(X"00");
	mem(152) := To_stdlogicvector(X"D1");
	mem(153) := To_stdlogicvector(X"BA");
	mem(154) := To_stdlogicvector(X"D2");
	mem(155) := To_stdlogicvector(X"BA");
	mem(156) := To_stdlogicvector(X"D3");
	mem(157) := To_stdlogicvector(X"BA");
	mem(158) := To_stdlogicvector(X"D4");
	mem(159) := To_stdlogicvector(X"BA");
	mem(160) := To_stdlogicvector(X"D5");
	mem(161) := To_stdlogicvector(X"BA");
	mem(162) := To_stdlogicvector(X"20");
	mem(163) := To_stdlogicvector(X"12");
	mem(164) := To_stdlogicvector(X"00");
	mem(165) := To_stdlogicvector(X"00");
	mem(166) := To_stdlogicvector(X"00");
	mem(167) := To_stdlogicvector(X"00");
	mem(168) := To_stdlogicvector(X"00");
	mem(169) := To_stdlogicvector(X"00");
	mem(170) := To_stdlogicvector(X"00");
	mem(171) := To_stdlogicvector(X"00");
	mem(172) := To_stdlogicvector(X"00");
	mem(173) := To_stdlogicvector(X"00");
	mem(174) := To_stdlogicvector(X"0A");
	mem(175) := To_stdlogicvector(X"0C");
	mem(176) := To_stdlogicvector(X"00");
	mem(177) := To_stdlogicvector(X"00");
	mem(178) := To_stdlogicvector(X"00");
	mem(179) := To_stdlogicvector(X"00");
	mem(180) := To_stdlogicvector(X"00");
	mem(181) := To_stdlogicvector(X"00");
	mem(182) := To_stdlogicvector(X"00");
	mem(183) := To_stdlogicvector(X"00");
	mem(184) := To_stdlogicvector(X"00");
	mem(185) := To_stdlogicvector(X"00");
	mem(186) := To_stdlogicvector(X"D1");
	mem(187) := To_stdlogicvector(X"BA");
	mem(188) := To_stdlogicvector(X"D2");
	mem(189) := To_stdlogicvector(X"BA");
	mem(190) := To_stdlogicvector(X"D3");
	mem(191) := To_stdlogicvector(X"BA");
	mem(192) := To_stdlogicvector(X"D4");
	mem(193) := To_stdlogicvector(X"BA");
	mem(194) := To_stdlogicvector(X"D5");
	mem(195) := To_stdlogicvector(X"BA");
	mem(196) := To_stdlogicvector(X"32");
	mem(197) := To_stdlogicvector(X"12");
	mem(198) := To_stdlogicvector(X"00");
	mem(199) := To_stdlogicvector(X"00");
	mem(200) := To_stdlogicvector(X"00");
	mem(201) := To_stdlogicvector(X"00");
	mem(202) := To_stdlogicvector(X"00");
	mem(203) := To_stdlogicvector(X"00");
	mem(204) := To_stdlogicvector(X"00");
	mem(205) := To_stdlogicvector(X"00");
	mem(206) := To_stdlogicvector(X"00");
	mem(207) := To_stdlogicvector(X"00");
	mem(208) := To_stdlogicvector(X"0A");
	mem(209) := To_stdlogicvector(X"0A");
	mem(210) := To_stdlogicvector(X"00");
	mem(211) := To_stdlogicvector(X"00");
	mem(212) := To_stdlogicvector(X"00");
	mem(213) := To_stdlogicvector(X"00");
	mem(214) := To_stdlogicvector(X"00");
	mem(215) := To_stdlogicvector(X"00");
	mem(216) := To_stdlogicvector(X"00");
	mem(217) := To_stdlogicvector(X"00");
	mem(218) := To_stdlogicvector(X"00");
	mem(219) := To_stdlogicvector(X"00");
	mem(220) := To_stdlogicvector(X"D1");
	mem(221) := To_stdlogicvector(X"BA");
	mem(222) := To_stdlogicvector(X"D2");
	mem(223) := To_stdlogicvector(X"BA");
	mem(224) := To_stdlogicvector(X"D3");
	mem(225) := To_stdlogicvector(X"BA");
	mem(226) := To_stdlogicvector(X"D4");
	mem(227) := To_stdlogicvector(X"BA");
	mem(228) := To_stdlogicvector(X"D5");
	mem(229) := To_stdlogicvector(X"BA");
	mem(230) := To_stdlogicvector(X"29");
	mem(231) := To_stdlogicvector(X"12");
	mem(232) := To_stdlogicvector(X"00");
	mem(233) := To_stdlogicvector(X"00");
	mem(234) := To_stdlogicvector(X"00");
	mem(235) := To_stdlogicvector(X"00");
	mem(236) := To_stdlogicvector(X"00");
	mem(237) := To_stdlogicvector(X"00");
	mem(238) := To_stdlogicvector(X"00");
	mem(239) := To_stdlogicvector(X"00");
	mem(240) := To_stdlogicvector(X"00");
	mem(241) := To_stdlogicvector(X"00");
	mem(242) := To_stdlogicvector(X"0A");
	mem(243) := To_stdlogicvector(X"0A");
	mem(244) := To_stdlogicvector(X"00");
	mem(245) := To_stdlogicvector(X"00");
	mem(246) := To_stdlogicvector(X"00");
	mem(247) := To_stdlogicvector(X"00");
	mem(248) := To_stdlogicvector(X"00");
	mem(249) := To_stdlogicvector(X"00");
	mem(250) := To_stdlogicvector(X"00");
	mem(251) := To_stdlogicvector(X"00");
	mem(252) := To_stdlogicvector(X"00");
	mem(253) := To_stdlogicvector(X"00");
	mem(254) := To_stdlogicvector(X"D1");
	mem(255) := To_stdlogicvector(X"BA");
	mem(256) := To_stdlogicvector(X"D2");
	mem(257) := To_stdlogicvector(X"BA");
	mem(258) := To_stdlogicvector(X"D3");
	mem(259) := To_stdlogicvector(X"BA");
	mem(260) := To_stdlogicvector(X"D4");
	mem(261) := To_stdlogicvector(X"BA");
	mem(262) := To_stdlogicvector(X"D5");
	mem(263) := To_stdlogicvector(X"BA");
	mem(264) := To_stdlogicvector(X"20");
	mem(265) := To_stdlogicvector(X"12");
	mem(266) := To_stdlogicvector(X"00");
	mem(267) := To_stdlogicvector(X"00");
	mem(268) := To_stdlogicvector(X"00");
	mem(269) := To_stdlogicvector(X"00");
	mem(270) := To_stdlogicvector(X"00");
	mem(271) := To_stdlogicvector(X"00");
	mem(272) := To_stdlogicvector(X"00");
	mem(273) := To_stdlogicvector(X"00");
	mem(274) := To_stdlogicvector(X"00");
	mem(275) := To_stdlogicvector(X"00");
	mem(276) := To_stdlogicvector(X"0A");
	mem(277) := To_stdlogicvector(X"06");
	mem(278) := To_stdlogicvector(X"00");
	mem(279) := To_stdlogicvector(X"00");
	mem(280) := To_stdlogicvector(X"00");
	mem(281) := To_stdlogicvector(X"00");
	mem(282) := To_stdlogicvector(X"00");
	mem(283) := To_stdlogicvector(X"00");
	mem(284) := To_stdlogicvector(X"00");
	mem(285) := To_stdlogicvector(X"00");
	mem(286) := To_stdlogicvector(X"00");
	mem(287) := To_stdlogicvector(X"00");
	mem(288) := To_stdlogicvector(X"D1");
	mem(289) := To_stdlogicvector(X"BA");
	mem(290) := To_stdlogicvector(X"D2");
	mem(291) := To_stdlogicvector(X"BA");
	mem(292) := To_stdlogicvector(X"D3");
	mem(293) := To_stdlogicvector(X"BA");
	mem(294) := To_stdlogicvector(X"D4");
	mem(295) := To_stdlogicvector(X"BA");
	mem(296) := To_stdlogicvector(X"D5");
	mem(297) := To_stdlogicvector(X"BA");
	mem(298) := To_stdlogicvector(X"2B");
	mem(299) := To_stdlogicvector(X"12");
	mem(300) := To_stdlogicvector(X"00");
	mem(301) := To_stdlogicvector(X"00");
	mem(302) := To_stdlogicvector(X"00");
	mem(303) := To_stdlogicvector(X"00");
	mem(304) := To_stdlogicvector(X"00");
	mem(305) := To_stdlogicvector(X"00");
	mem(306) := To_stdlogicvector(X"00");
	mem(307) := To_stdlogicvector(X"00");
	mem(308) := To_stdlogicvector(X"00");
	mem(309) := To_stdlogicvector(X"00");
	mem(310) := To_stdlogicvector(X"0A");
	mem(311) := To_stdlogicvector(X"06");
	mem(312) := To_stdlogicvector(X"00");
	mem(313) := To_stdlogicvector(X"00");
	mem(314) := To_stdlogicvector(X"00");
	mem(315) := To_stdlogicvector(X"00");
	mem(316) := To_stdlogicvector(X"00");
	mem(317) := To_stdlogicvector(X"00");
	mem(318) := To_stdlogicvector(X"00");
	mem(319) := To_stdlogicvector(X"00");
	mem(320) := To_stdlogicvector(X"00");
	mem(321) := To_stdlogicvector(X"00");
	mem(322) := To_stdlogicvector(X"D1");
	mem(323) := To_stdlogicvector(X"BA");
	mem(324) := To_stdlogicvector(X"D2");
	mem(325) := To_stdlogicvector(X"BA");
	mem(326) := To_stdlogicvector(X"D3");
	mem(327) := To_stdlogicvector(X"BA");
	mem(328) := To_stdlogicvector(X"D4");
	mem(329) := To_stdlogicvector(X"BA");
	mem(330) := To_stdlogicvector(X"D5");
	mem(331) := To_stdlogicvector(X"BA");
	mem(332) := To_stdlogicvector(X"00");
	mem(333) := To_stdlogicvector(X"00");
	mem(334) := To_stdlogicvector(X"00");
	mem(335) := To_stdlogicvector(X"00");
	mem(336) := To_stdlogicvector(X"00");
	mem(337) := To_stdlogicvector(X"00");
	mem(338) := To_stdlogicvector(X"00");
	mem(339) := To_stdlogicvector(X"00");
	mem(340) := To_stdlogicvector(X"00");
	mem(341) := To_stdlogicvector(X"00");
	mem(342) := To_stdlogicvector(X"FA");
	mem(343) := To_stdlogicvector(X"0F");
	mem(344) := To_stdlogicvector(X"00");
	mem(345) := To_stdlogicvector(X"00");
	mem(346) := To_stdlogicvector(X"00");
	mem(347) := To_stdlogicvector(X"00");
	mem(348) := To_stdlogicvector(X"00");
	mem(349) := To_stdlogicvector(X"00");
	mem(350) := To_stdlogicvector(X"00");
	mem(351) := To_stdlogicvector(X"00");
	mem(352) := To_stdlogicvector(X"00");
	mem(353) := To_stdlogicvector(X"00");
	mem(354) := To_stdlogicvector(X"DD");
	mem(355) := To_stdlogicvector(X"BA");
