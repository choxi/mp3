	mem(0) := To_stdlogicvector(X"0A");
	mem(1) := To_stdlogicvector(X"F0");
	mem(2) := To_stdlogicvector(X"13");
	mem(3) := To_stdlogicvector(X"E2");
	mem(4) := To_stdlogicvector(X"40");
	mem(5) := To_stdlogicvector(X"C0");
	mem(6) := To_stdlogicvector(X"21");
	mem(7) := To_stdlogicvector(X"10");
	mem(8) := To_stdlogicvector(X"21");
	mem(9) := To_stdlogicvector(X"10");
	mem(10) := To_stdlogicvector(X"21");
	mem(11) := To_stdlogicvector(X"10");
	mem(12) := To_stdlogicvector(X"21");
	mem(13) := To_stdlogicvector(X"10");
	mem(14) := To_stdlogicvector(X"21");
	mem(15) := To_stdlogicvector(X"10");
	mem(16) := To_stdlogicvector(X"21");
	mem(17) := To_stdlogicvector(X"10");
	mem(18) := To_stdlogicvector(X"21");
	mem(19) := To_stdlogicvector(X"10");
	mem(20) := To_stdlogicvector(X"26");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"21");
	mem(23) := To_stdlogicvector(X"10");
	mem(24) := To_stdlogicvector(X"21");
	mem(25) := To_stdlogicvector(X"10");
	mem(26) := To_stdlogicvector(X"21");
	mem(27) := To_stdlogicvector(X"10");
	mem(28) := To_stdlogicvector(X"21");
	mem(29) := To_stdlogicvector(X"10");
	mem(30) := To_stdlogicvector(X"21");
	mem(31) := To_stdlogicvector(X"10");
	mem(32) := To_stdlogicvector(X"21");
	mem(33) := To_stdlogicvector(X"10");
	mem(34) := To_stdlogicvector(X"21");
	mem(35) := To_stdlogicvector(X"10");
	mem(36) := To_stdlogicvector(X"21");
	mem(37) := To_stdlogicvector(X"10");
	mem(38) := To_stdlogicvector(X"2F");
	mem(39) := To_stdlogicvector(X"19");
	mem(40) := To_stdlogicvector(X"C0");
	mem(41) := To_stdlogicvector(X"C1");
	mem(42) := To_stdlogicvector(X"FF");
	mem(43) := To_stdlogicvector(X"0F");
