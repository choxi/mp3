	mem(0) := To_stdlogicvector(X"FF");
	mem(1) := To_stdlogicvector(X"E1");
	mem(2) := To_stdlogicvector(X"20");
	mem(3) := To_stdlogicvector(X"52");
	mem(4) := To_stdlogicvector(X"20");
	mem(5) := To_stdlogicvector(X"54");
	mem(6) := To_stdlogicvector(X"20");
	mem(7) := To_stdlogicvector(X"56");
	mem(8) := To_stdlogicvector(X"20");
	mem(9) := To_stdlogicvector(X"58");
	mem(10) := To_stdlogicvector(X"20");
	mem(11) := To_stdlogicvector(X"5A");
	mem(12) := To_stdlogicvector(X"A0");
	mem(13) := To_stdlogicvector(X"5D");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"22");
	mem(17) := To_stdlogicvector(X"10");
	mem(18) := To_stdlogicvector(X"10");
	mem(19) := To_stdlogicvector(X"A2");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"00");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"00");
	mem(25) := To_stdlogicvector(X"00");
	mem(26) := To_stdlogicvector(X"00");
	mem(27) := To_stdlogicvector(X"00");
	mem(28) := To_stdlogicvector(X"00");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"10");
	mem(31) := To_stdlogicvector(X"0E");
	mem(32) := To_stdlogicvector(X"DD");
	mem(33) := To_stdlogicvector(X"BA");
	mem(34) := To_stdlogicvector(X"30");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"DD");
	mem(37) := To_stdlogicvector(X"BA");
	mem(38) := To_stdlogicvector(X"DD");
	mem(39) := To_stdlogicvector(X"BA");
	mem(40) := To_stdlogicvector(X"DD");
	mem(41) := To_stdlogicvector(X"BA");
	mem(42) := To_stdlogicvector(X"DD");
	mem(43) := To_stdlogicvector(X"BA");
	mem(44) := To_stdlogicvector(X"DD");
	mem(45) := To_stdlogicvector(X"BA");
	mem(46) := To_stdlogicvector(X"DD");
	mem(47) := To_stdlogicvector(X"BA");
	mem(48) := To_stdlogicvector(X"0D");
	mem(49) := To_stdlogicvector(X"60");
	mem(50) := To_stdlogicvector(X"DD");
	mem(51) := To_stdlogicvector(X"BA");
	mem(52) := To_stdlogicvector(X"DD");
	mem(53) := To_stdlogicvector(X"BA");
	mem(54) := To_stdlogicvector(X"DD");
	mem(55) := To_stdlogicvector(X"BA");
	mem(56) := To_stdlogicvector(X"DD");
	mem(57) := To_stdlogicvector(X"BA");
	mem(58) := To_stdlogicvector(X"DD");
	mem(59) := To_stdlogicvector(X"BA");
	mem(60) := To_stdlogicvector(X"DD");
	mem(61) := To_stdlogicvector(X"BA");
	mem(62) := To_stdlogicvector(X"DD");
	mem(63) := To_stdlogicvector(X"BA");
	mem(64) := To_stdlogicvector(X"FF");
	mem(65) := To_stdlogicvector(X"E1");
	mem(66) := To_stdlogicvector(X"20");
	mem(67) := To_stdlogicvector(X"52");
	mem(68) := To_stdlogicvector(X"20");
	mem(69) := To_stdlogicvector(X"54");
	mem(70) := To_stdlogicvector(X"20");
	mem(71) := To_stdlogicvector(X"56");
	mem(72) := To_stdlogicvector(X"20");
	mem(73) := To_stdlogicvector(X"58");
	mem(74) := To_stdlogicvector(X"20");
	mem(75) := To_stdlogicvector(X"5A");
	mem(76) := To_stdlogicvector(X"A1");
	mem(77) := To_stdlogicvector(X"1D");
	mem(78) := To_stdlogicvector(X"00");
	mem(79) := To_stdlogicvector(X"00");
	mem(80) := To_stdlogicvector(X"90");
	mem(81) := To_stdlogicvector(X"64");
	mem(82) := To_stdlogicvector(X"22");
	mem(83) := To_stdlogicvector(X"10");
	mem(84) := To_stdlogicvector(X"10");
	mem(85) := To_stdlogicvector(X"A2");
	mem(86) := To_stdlogicvector(X"00");
	mem(87) := To_stdlogicvector(X"00");
	mem(88) := To_stdlogicvector(X"00");
	mem(89) := To_stdlogicvector(X"00");
	mem(90) := To_stdlogicvector(X"00");
	mem(91) := To_stdlogicvector(X"00");
	mem(92) := To_stdlogicvector(X"00");
	mem(93) := To_stdlogicvector(X"00");
	mem(94) := To_stdlogicvector(X"10");
	mem(95) := To_stdlogicvector(X"0E");
	mem(96) := To_stdlogicvector(X"DD");
	mem(97) := To_stdlogicvector(X"BA");
	mem(98) := To_stdlogicvector(X"70");
	mem(99) := To_stdlogicvector(X"00");
	mem(100) := To_stdlogicvector(X"DD");
	mem(101) := To_stdlogicvector(X"BA");
	mem(102) := To_stdlogicvector(X"DD");
	mem(103) := To_stdlogicvector(X"BA");
	mem(104) := To_stdlogicvector(X"DD");
	mem(105) := To_stdlogicvector(X"BA");
	mem(106) := To_stdlogicvector(X"DD");
	mem(107) := To_stdlogicvector(X"BA");
	mem(108) := To_stdlogicvector(X"DD");
	mem(109) := To_stdlogicvector(X"BA");
	mem(110) := To_stdlogicvector(X"DD");
	mem(111) := To_stdlogicvector(X"BA");
	mem(112) := To_stdlogicvector(X"0D");
	mem(113) := To_stdlogicvector(X"60");
	mem(114) := To_stdlogicvector(X"DD");
	mem(115) := To_stdlogicvector(X"BA");
	mem(116) := To_stdlogicvector(X"DD");
	mem(117) := To_stdlogicvector(X"BA");
	mem(118) := To_stdlogicvector(X"DD");
	mem(119) := To_stdlogicvector(X"BA");
	mem(120) := To_stdlogicvector(X"DD");
	mem(121) := To_stdlogicvector(X"BA");
	mem(122) := To_stdlogicvector(X"DD");
	mem(123) := To_stdlogicvector(X"BA");
	mem(124) := To_stdlogicvector(X"DD");
	mem(125) := To_stdlogicvector(X"BA");
	mem(126) := To_stdlogicvector(X"DD");
	mem(127) := To_stdlogicvector(X"BA");
	mem(128) := To_stdlogicvector(X"FF");
	mem(129) := To_stdlogicvector(X"E1");
	mem(130) := To_stdlogicvector(X"20");
	mem(131) := To_stdlogicvector(X"52");
	mem(132) := To_stdlogicvector(X"20");
	mem(133) := To_stdlogicvector(X"54");
	mem(134) := To_stdlogicvector(X"20");
	mem(135) := To_stdlogicvector(X"56");
	mem(136) := To_stdlogicvector(X"20");
	mem(137) := To_stdlogicvector(X"58");
	mem(138) := To_stdlogicvector(X"20");
	mem(139) := To_stdlogicvector(X"5A");
	mem(140) := To_stdlogicvector(X"A1");
	mem(141) := To_stdlogicvector(X"1D");
	mem(142) := To_stdlogicvector(X"00");
	mem(143) := To_stdlogicvector(X"00");
	mem(144) := To_stdlogicvector(X"10");
	mem(145) := To_stdlogicvector(X"64");
	mem(146) := To_stdlogicvector(X"22");
	mem(147) := To_stdlogicvector(X"10");
	mem(148) := To_stdlogicvector(X"10");
	mem(149) := To_stdlogicvector(X"A2");
	mem(150) := To_stdlogicvector(X"00");
	mem(151) := To_stdlogicvector(X"00");
	mem(152) := To_stdlogicvector(X"00");
	mem(153) := To_stdlogicvector(X"00");
	mem(154) := To_stdlogicvector(X"00");
	mem(155) := To_stdlogicvector(X"00");
	mem(156) := To_stdlogicvector(X"00");
	mem(157) := To_stdlogicvector(X"00");
	mem(158) := To_stdlogicvector(X"08");
	mem(159) := To_stdlogicvector(X"0E");
	mem(160) := To_stdlogicvector(X"0D");
	mem(161) := To_stdlogicvector(X"60");
	mem(162) := To_stdlogicvector(X"A8");
	mem(163) := To_stdlogicvector(X"00");
	mem(164) := To_stdlogicvector(X"DD");
	mem(165) := To_stdlogicvector(X"BA");
	mem(166) := To_stdlogicvector(X"DD");
	mem(167) := To_stdlogicvector(X"BA");
	mem(168) := To_stdlogicvector(X"0D");
	mem(169) := To_stdlogicvector(X"60");
	mem(170) := To_stdlogicvector(X"DD");
	mem(171) := To_stdlogicvector(X"BA");
	mem(172) := To_stdlogicvector(X"DD");
	mem(173) := To_stdlogicvector(X"BA");
	mem(174) := To_stdlogicvector(X"DD");
	mem(175) := To_stdlogicvector(X"BA");
	mem(176) := To_stdlogicvector(X"FF");
	mem(177) := To_stdlogicvector(X"E1");
	mem(178) := To_stdlogicvector(X"20");
	mem(179) := To_stdlogicvector(X"52");
	mem(180) := To_stdlogicvector(X"20");
	mem(181) := To_stdlogicvector(X"54");
	mem(182) := To_stdlogicvector(X"20");
	mem(183) := To_stdlogicvector(X"56");
	mem(184) := To_stdlogicvector(X"20");
	mem(185) := To_stdlogicvector(X"58");
	mem(186) := To_stdlogicvector(X"20");
	mem(187) := To_stdlogicvector(X"5A");
	mem(188) := To_stdlogicvector(X"A1");
	mem(189) := To_stdlogicvector(X"1D");
	mem(190) := To_stdlogicvector(X"00");
	mem(191) := To_stdlogicvector(X"00");
	mem(192) := To_stdlogicvector(X"22");
	mem(193) := To_stdlogicvector(X"10");
	mem(194) := To_stdlogicvector(X"10");
	mem(195) := To_stdlogicvector(X"A2");
	mem(196) := To_stdlogicvector(X"00");
	mem(197) := To_stdlogicvector(X"00");
	mem(198) := To_stdlogicvector(X"00");
	mem(199) := To_stdlogicvector(X"00");
	mem(200) := To_stdlogicvector(X"00");
	mem(201) := To_stdlogicvector(X"00");
	mem(202) := To_stdlogicvector(X"00");
	mem(203) := To_stdlogicvector(X"00");
	mem(204) := To_stdlogicvector(X"00");
	mem(205) := To_stdlogicvector(X"00");
	mem(206) := To_stdlogicvector(X"08");
	mem(207) := To_stdlogicvector(X"0E");
	mem(208) := To_stdlogicvector(X"DD");
	mem(209) := To_stdlogicvector(X"BA");
	mem(210) := To_stdlogicvector(X"D8");
	mem(211) := To_stdlogicvector(X"00");
	mem(212) := To_stdlogicvector(X"DD");
	mem(213) := To_stdlogicvector(X"BA");
	mem(214) := To_stdlogicvector(X"DD");
	mem(215) := To_stdlogicvector(X"BA");
	mem(216) := To_stdlogicvector(X"0D");
	mem(217) := To_stdlogicvector(X"60");
	mem(218) := To_stdlogicvector(X"DD");
	mem(219) := To_stdlogicvector(X"BA");
	mem(220) := To_stdlogicvector(X"DD");
	mem(221) := To_stdlogicvector(X"BA");
	mem(222) := To_stdlogicvector(X"DD");
	mem(223) := To_stdlogicvector(X"BA");
	mem(224) := To_stdlogicvector(X"20");
	mem(225) := To_stdlogicvector(X"50");
	mem(226) := To_stdlogicvector(X"20");
	mem(227) := To_stdlogicvector(X"52");
	mem(228) := To_stdlogicvector(X"20");
	mem(229) := To_stdlogicvector(X"54");
	mem(230) := To_stdlogicvector(X"20");
	mem(231) := To_stdlogicvector(X"56");
	mem(232) := To_stdlogicvector(X"20");
	mem(233) := To_stdlogicvector(X"58");
	mem(234) := To_stdlogicvector(X"20");
	mem(235) := To_stdlogicvector(X"5A");
	mem(236) := To_stdlogicvector(X"A1");
	mem(237) := To_stdlogicvector(X"1D");
	mem(238) := To_stdlogicvector(X"00");
	mem(239) := To_stdlogicvector(X"00");
	mem(240) := To_stdlogicvector(X"02");
	mem(241) := To_stdlogicvector(X"E4");
	mem(242) := To_stdlogicvector(X"80");
	mem(243) := To_stdlogicvector(X"C0");
	mem(244) := To_stdlogicvector(X"02");
	mem(245) := To_stdlogicvector(X"0E");
	mem(246) := To_stdlogicvector(X"66");
	mem(247) := To_stdlogicvector(X"12");
	mem(248) := To_stdlogicvector(X"03");
	mem(249) := To_stdlogicvector(X"0E");
	mem(250) := To_stdlogicvector(X"65");
	mem(251) := To_stdlogicvector(X"12");
	mem(252) := To_stdlogicvector(X"00");
	mem(253) := To_stdlogicvector(X"00");
	mem(254) := To_stdlogicvector(X"00");
	mem(255) := To_stdlogicvector(X"0E");
	mem(256) := To_stdlogicvector(X"FF");
	mem(257) := To_stdlogicvector(X"E1");
	mem(258) := To_stdlogicvector(X"20");
	mem(259) := To_stdlogicvector(X"52");
	mem(260) := To_stdlogicvector(X"20");
	mem(261) := To_stdlogicvector(X"54");
	mem(262) := To_stdlogicvector(X"20");
	mem(263) := To_stdlogicvector(X"56");
	mem(264) := To_stdlogicvector(X"20");
	mem(265) := To_stdlogicvector(X"58");
	mem(266) := To_stdlogicvector(X"20");
	mem(267) := To_stdlogicvector(X"5A");
	mem(268) := To_stdlogicvector(X"A1");
	mem(269) := To_stdlogicvector(X"1D");
	mem(270) := To_stdlogicvector(X"00");
	mem(271) := To_stdlogicvector(X"00");
	mem(272) := To_stdlogicvector(X"10");
	mem(273) := To_stdlogicvector(X"64");
	mem(274) := To_stdlogicvector(X"80");
	mem(275) := To_stdlogicvector(X"C0");
	mem(276) := To_stdlogicvector(X"0A");
	mem(277) := To_stdlogicvector(X"0E");
	mem(278) := To_stdlogicvector(X"00");
	mem(279) := To_stdlogicvector(X"00");
	mem(280) := To_stdlogicvector(X"00");
	mem(281) := To_stdlogicvector(X"00");
	mem(282) := To_stdlogicvector(X"00");
	mem(283) := To_stdlogicvector(X"00");
	mem(284) := To_stdlogicvector(X"00");
	mem(285) := To_stdlogicvector(X"00");
	mem(286) := To_stdlogicvector(X"00");
	mem(287) := To_stdlogicvector(X"00");
	mem(288) := To_stdlogicvector(X"26");
	mem(289) := To_stdlogicvector(X"01");
	mem(290) := To_stdlogicvector(X"00");
	mem(291) := To_stdlogicvector(X"00");
	mem(292) := To_stdlogicvector(X"00");
	mem(293) := To_stdlogicvector(X"00");
	mem(294) := To_stdlogicvector(X"66");
	mem(295) := To_stdlogicvector(X"12");
	mem(296) := To_stdlogicvector(X"03");
	mem(297) := To_stdlogicvector(X"0E");
	mem(298) := To_stdlogicvector(X"65");
	mem(299) := To_stdlogicvector(X"12");
	mem(300) := To_stdlogicvector(X"01");
	mem(301) := To_stdlogicvector(X"0E");
	mem(302) := To_stdlogicvector(X"00");
	mem(303) := To_stdlogicvector(X"00");
	mem(304) := To_stdlogicvector(X"20");
	mem(305) := To_stdlogicvector(X"50");
	mem(306) := To_stdlogicvector(X"20");
	mem(307) := To_stdlogicvector(X"52");
	mem(308) := To_stdlogicvector(X"20");
	mem(309) := To_stdlogicvector(X"54");
	mem(310) := To_stdlogicvector(X"20");
	mem(311) := To_stdlogicvector(X"56");
	mem(312) := To_stdlogicvector(X"20");
	mem(313) := To_stdlogicvector(X"58");
	mem(314) := To_stdlogicvector(X"20");
	mem(315) := To_stdlogicvector(X"5A");
	mem(316) := To_stdlogicvector(X"A1");
	mem(317) := To_stdlogicvector(X"1D");
	mem(318) := To_stdlogicvector(X"00");
	mem(319) := To_stdlogicvector(X"00");
	mem(320) := To_stdlogicvector(X"03");
	mem(321) := To_stdlogicvector(X"EE");
	mem(322) := To_stdlogicvector(X"C0");
	mem(323) := To_stdlogicvector(X"C1");
	mem(324) := To_stdlogicvector(X"03");
	mem(325) := To_stdlogicvector(X"0E");
	mem(326) := To_stdlogicvector(X"00");
	mem(327) := To_stdlogicvector(X"00");
	mem(328) := To_stdlogicvector(X"66");
	mem(329) := To_stdlogicvector(X"12");
	mem(330) := To_stdlogicvector(X"02");
	mem(331) := To_stdlogicvector(X"0E");
	mem(332) := To_stdlogicvector(X"65");
	mem(333) := To_stdlogicvector(X"12");
	mem(334) := To_stdlogicvector(X"00");
	mem(335) := To_stdlogicvector(X"0E");
	mem(336) := To_stdlogicvector(X"20");
	mem(337) := To_stdlogicvector(X"50");
	mem(338) := To_stdlogicvector(X"20");
	mem(339) := To_stdlogicvector(X"52");
	mem(340) := To_stdlogicvector(X"20");
	mem(341) := To_stdlogicvector(X"54");
	mem(342) := To_stdlogicvector(X"20");
	mem(343) := To_stdlogicvector(X"56");
	mem(344) := To_stdlogicvector(X"20");
	mem(345) := To_stdlogicvector(X"58");
	mem(346) := To_stdlogicvector(X"20");
	mem(347) := To_stdlogicvector(X"5A");
	mem(348) := To_stdlogicvector(X"A1");
	mem(349) := To_stdlogicvector(X"1D");
	mem(350) := To_stdlogicvector(X"00");
	mem(351) := To_stdlogicvector(X"00");
	mem(352) := To_stdlogicvector(X"0A");
	mem(353) := To_stdlogicvector(X"E4");
	mem(354) := To_stdlogicvector(X"80");
	mem(355) := To_stdlogicvector(X"40");
	mem(356) := To_stdlogicvector(X"0A");
	mem(357) := To_stdlogicvector(X"0E");
	mem(358) := To_stdlogicvector(X"66");
	mem(359) := To_stdlogicvector(X"12");
	mem(360) := To_stdlogicvector(X"0B");
	mem(361) := To_stdlogicvector(X"0E");
	mem(362) := To_stdlogicvector(X"07");
	mem(363) := To_stdlogicvector(X"0E");
	mem(364) := To_stdlogicvector(X"06");
	mem(365) := To_stdlogicvector(X"0E");
	mem(366) := To_stdlogicvector(X"05");
	mem(367) := To_stdlogicvector(X"0E");
	mem(368) := To_stdlogicvector(X"00");
	mem(369) := To_stdlogicvector(X"00");
	mem(370) := To_stdlogicvector(X"00");
	mem(371) := To_stdlogicvector(X"00");
	mem(372) := To_stdlogicvector(X"00");
	mem(373) := To_stdlogicvector(X"00");
	mem(374) := To_stdlogicvector(X"E2");
	mem(375) := To_stdlogicvector(X"1F");
	mem(376) := To_stdlogicvector(X"C0");
	mem(377) := To_stdlogicvector(X"C1");
	mem(378) := To_stdlogicvector(X"65");
	mem(379) := To_stdlogicvector(X"12");
	mem(380) := To_stdlogicvector(X"01");
	mem(381) := To_stdlogicvector(X"0E");
	mem(382) := To_stdlogicvector(X"00");
	mem(383) := To_stdlogicvector(X"00");
	mem(384) := To_stdlogicvector(X"FF");
	mem(385) := To_stdlogicvector(X"E1");
	mem(386) := To_stdlogicvector(X"20");
	mem(387) := To_stdlogicvector(X"52");
	mem(388) := To_stdlogicvector(X"20");
	mem(389) := To_stdlogicvector(X"54");
	mem(390) := To_stdlogicvector(X"20");
	mem(391) := To_stdlogicvector(X"56");
	mem(392) := To_stdlogicvector(X"20");
	mem(393) := To_stdlogicvector(X"58");
	mem(394) := To_stdlogicvector(X"20");
	mem(395) := To_stdlogicvector(X"5A");
	mem(396) := To_stdlogicvector(X"A1");
	mem(397) := To_stdlogicvector(X"1D");
	mem(398) := To_stdlogicvector(X"E0");
	mem(399) := To_stdlogicvector(X"5F");
	mem(400) := To_stdlogicvector(X"E6");
	mem(401) := To_stdlogicvector(X"16");
	mem(402) := To_stdlogicvector(X"11");
	mem(403) := To_stdlogicvector(X"64");
	mem(404) := To_stdlogicvector(X"80");
	mem(405) := To_stdlogicvector(X"76");
	mem(406) := To_stdlogicvector(X"00");
	mem(407) := To_stdlogicvector(X"00");
	mem(408) := To_stdlogicvector(X"80");
	mem(409) := To_stdlogicvector(X"62");
	mem(410) := To_stdlogicvector(X"00");
	mem(411) := To_stdlogicvector(X"00");
	mem(412) := To_stdlogicvector(X"00");
	mem(413) := To_stdlogicvector(X"00");
	mem(414) := To_stdlogicvector(X"08");
	mem(415) := To_stdlogicvector(X"0E");
	mem(416) := To_stdlogicvector(X"DD");
	mem(417) := To_stdlogicvector(X"BA");
	mem(418) := To_stdlogicvector(X"A8");
	mem(419) := To_stdlogicvector(X"01");
	mem(420) := To_stdlogicvector(X"DD");
	mem(421) := To_stdlogicvector(X"BA");
	mem(422) := To_stdlogicvector(X"DD");
	mem(423) := To_stdlogicvector(X"BA");
	mem(424) := To_stdlogicvector(X"DD");
	mem(425) := To_stdlogicvector(X"BA");
	mem(426) := To_stdlogicvector(X"DD");
	mem(427) := To_stdlogicvector(X"BA");
	mem(428) := To_stdlogicvector(X"DD");
	mem(429) := To_stdlogicvector(X"BA");
	mem(430) := To_stdlogicvector(X"DD");
	mem(431) := To_stdlogicvector(X"BA");
	mem(432) := To_stdlogicvector(X"FF");
	mem(433) := To_stdlogicvector(X"0F");
