	mem(0) := To_stdlogicvector(X"F9");
	mem(1) := To_stdlogicvector(X"E0");
	mem(2) := To_stdlogicvector(X"6C");
	mem(3) := To_stdlogicvector(X"12");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"7B");
	mem(11) := To_stdlogicvector(X"12");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"00");
	mem(14) := To_stdlogicvector(X"00");
	mem(15) := To_stdlogicvector(X"00");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"60");
	mem(19) := To_stdlogicvector(X"12");
	mem(20) := To_stdlogicvector(X"00");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"00");
	mem(23) := To_stdlogicvector(X"00");
	mem(24) := To_stdlogicvector(X"00");
	mem(25) := To_stdlogicvector(X"00");
	mem(26) := To_stdlogicvector(X"10");
	mem(27) := To_stdlogicvector(X"72");
	mem(28) := To_stdlogicvector(X"2F");
	mem(29) := To_stdlogicvector(X"54");
	mem(30) := To_stdlogicvector(X"00");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"00");
	mem(33) := To_stdlogicvector(X"00");
	mem(34) := To_stdlogicvector(X"00");
	mem(35) := To_stdlogicvector(X"00");
	mem(36) := To_stdlogicvector(X"11");
	mem(37) := To_stdlogicvector(X"74");
	mem(38) := To_stdlogicvector(X"00");
	mem(39) := To_stdlogicvector(X"00");
	mem(40) := To_stdlogicvector(X"00");
	mem(41) := To_stdlogicvector(X"00");
	mem(42) := To_stdlogicvector(X"00");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"04");
	mem(45) := To_stdlogicvector(X"66");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"00");
	mem(49) := To_stdlogicvector(X"00");
	mem(50) := To_stdlogicvector(X"00");
	mem(51) := To_stdlogicvector(X"00");
	mem(52) := To_stdlogicvector(X"05");
	mem(53) := To_stdlogicvector(X"68");
	mem(54) := To_stdlogicvector(X"00");
	mem(55) := To_stdlogicvector(X"00");
	mem(56) := To_stdlogicvector(X"00");
	mem(57) := To_stdlogicvector(X"00");
	mem(58) := To_stdlogicvector(X"00");
	mem(59) := To_stdlogicvector(X"00");
	mem(60) := To_stdlogicvector(X"06");
	mem(61) := To_stdlogicvector(X"6A");
	mem(62) := To_stdlogicvector(X"00");
	mem(63) := To_stdlogicvector(X"00");
	mem(64) := To_stdlogicvector(X"00");
	mem(65) := To_stdlogicvector(X"00");
	mem(66) := To_stdlogicvector(X"00");
	mem(67) := To_stdlogicvector(X"00");
	mem(68) := To_stdlogicvector(X"07");
	mem(69) := To_stdlogicvector(X"6C");
	mem(70) := To_stdlogicvector(X"00");
	mem(71) := To_stdlogicvector(X"00");
	mem(72) := To_stdlogicvector(X"00");
	mem(73) := To_stdlogicvector(X"00");
	mem(74) := To_stdlogicvector(X"00");
	mem(75) := To_stdlogicvector(X"00");
	mem(76) := To_stdlogicvector(X"C4");
	mem(77) := To_stdlogicvector(X"16");
	mem(78) := To_stdlogicvector(X"00");
	mem(79) := To_stdlogicvector(X"00");
	mem(80) := To_stdlogicvector(X"00");
	mem(81) := To_stdlogicvector(X"00");
	mem(82) := To_stdlogicvector(X"00");
	mem(83) := To_stdlogicvector(X"00");
	mem(84) := To_stdlogicvector(X"C3");
	mem(85) := To_stdlogicvector(X"16");
	mem(86) := To_stdlogicvector(X"00");
	mem(87) := To_stdlogicvector(X"00");
	mem(88) := To_stdlogicvector(X"00");
	mem(89) := To_stdlogicvector(X"00");
	mem(90) := To_stdlogicvector(X"00");
	mem(91) := To_stdlogicvector(X"00");
	mem(92) := To_stdlogicvector(X"12");
	mem(93) := To_stdlogicvector(X"76");
	mem(94) := To_stdlogicvector(X"43");
	mem(95) := To_stdlogicvector(X"59");
	mem(96) := To_stdlogicvector(X"00");
	mem(97) := To_stdlogicvector(X"00");
	mem(98) := To_stdlogicvector(X"00");
	mem(99) := To_stdlogicvector(X"00");
	mem(100) := To_stdlogicvector(X"00");
	mem(101) := To_stdlogicvector(X"00");
	mem(102) := To_stdlogicvector(X"11");
	mem(103) := To_stdlogicvector(X"78");
	mem(104) := To_stdlogicvector(X"7F");
	mem(105) := To_stdlogicvector(X"9B");
	mem(106) := To_stdlogicvector(X"00");
	mem(107) := To_stdlogicvector(X"00");
	mem(108) := To_stdlogicvector(X"00");
	mem(109) := To_stdlogicvector(X"00");
	mem(110) := To_stdlogicvector(X"00");
	mem(111) := To_stdlogicvector(X"00");
	mem(112) := To_stdlogicvector(X"14");
	mem(113) := To_stdlogicvector(X"7A");
	mem(114) := To_stdlogicvector(X"08");
	mem(115) := To_stdlogicvector(X"6C");
	mem(116) := To_stdlogicvector(X"00");
	mem(117) := To_stdlogicvector(X"00");
	mem(118) := To_stdlogicvector(X"00");
	mem(119) := To_stdlogicvector(X"00");
	mem(120) := To_stdlogicvector(X"00");
	mem(121) := To_stdlogicvector(X"00");
	mem(122) := To_stdlogicvector(X"08");
	mem(123) := To_stdlogicvector(X"6E");
	mem(124) := To_stdlogicvector(X"00");
	mem(125) := To_stdlogicvector(X"00");
	mem(126) := To_stdlogicvector(X"00");
	mem(127) := To_stdlogicvector(X"00");
	mem(128) := To_stdlogicvector(X"00");
	mem(129) := To_stdlogicvector(X"00");
	mem(130) := To_stdlogicvector(X"A8");
	mem(131) := To_stdlogicvector(X"DD");
	mem(132) := To_stdlogicvector(X"00");
	mem(133) := To_stdlogicvector(X"00");
	mem(134) := To_stdlogicvector(X"00");
	mem(135) := To_stdlogicvector(X"00");
	mem(136) := To_stdlogicvector(X"00");
	mem(137) := To_stdlogicvector(X"00");
	mem(138) := To_stdlogicvector(X"D3");
	mem(139) := To_stdlogicvector(X"DF");
	mem(140) := To_stdlogicvector(X"00");
	mem(141) := To_stdlogicvector(X"00");
	mem(142) := To_stdlogicvector(X"00");
	mem(143) := To_stdlogicvector(X"00");
	mem(144) := To_stdlogicvector(X"00");
	mem(145) := To_stdlogicvector(X"00");
	mem(146) := To_stdlogicvector(X"B6");
	mem(147) := To_stdlogicvector(X"DD");
	mem(148) := To_stdlogicvector(X"00");
	mem(149) := To_stdlogicvector(X"00");
	mem(150) := To_stdlogicvector(X"00");
	mem(151) := To_stdlogicvector(X"00");
	mem(152) := To_stdlogicvector(X"00");
	mem(153) := To_stdlogicvector(X"00");
	mem(154) := To_stdlogicvector(X"13");
	mem(155) := To_stdlogicvector(X"7C");
	mem(156) := To_stdlogicvector(X"00");
	mem(157) := To_stdlogicvector(X"00");
	mem(158) := To_stdlogicvector(X"00");
	mem(159) := To_stdlogicvector(X"00");
	mem(160) := To_stdlogicvector(X"00");
	mem(161) := To_stdlogicvector(X"00");
	mem(162) := To_stdlogicvector(X"13");
	mem(163) := To_stdlogicvector(X"7E");
	mem(164) := To_stdlogicvector(X"00");
	mem(165) := To_stdlogicvector(X"00");
	mem(166) := To_stdlogicvector(X"00");
	mem(167) := To_stdlogicvector(X"00");
	mem(168) := To_stdlogicvector(X"00");
	mem(169) := To_stdlogicvector(X"00");
	mem(170) := To_stdlogicvector(X"00");
	mem(171) := To_stdlogicvector(X"62");
	mem(172) := To_stdlogicvector(X"00");
	mem(173) := To_stdlogicvector(X"64");
	mem(174) := To_stdlogicvector(X"06");
	mem(175) := To_stdlogicvector(X"66");
	mem(176) := To_stdlogicvector(X"07");
	mem(177) := To_stdlogicvector(X"68");
	mem(178) := To_stdlogicvector(X"08");
	mem(179) := To_stdlogicvector(X"6A");
	mem(180) := To_stdlogicvector(X"04");
	mem(181) := To_stdlogicvector(X"6C");
	mem(182) := To_stdlogicvector(X"05");
	mem(183) := To_stdlogicvector(X"6E");
	mem(184) := To_stdlogicvector(X"09");
	mem(185) := To_stdlogicvector(X"62");
	mem(186) := To_stdlogicvector(X"00");
	mem(187) := To_stdlogicvector(X"00");
	mem(188) := To_stdlogicvector(X"00");
	mem(189) := To_stdlogicvector(X"00");
	mem(190) := To_stdlogicvector(X"00");
	mem(191) := To_stdlogicvector(X"00");
	mem(192) := To_stdlogicvector(X"0B");
	mem(193) := To_stdlogicvector(X"E4");
	mem(194) := To_stdlogicvector(X"00");
	mem(195) := To_stdlogicvector(X"00");
	mem(196) := To_stdlogicvector(X"00");
	mem(197) := To_stdlogicvector(X"00");
	mem(198) := To_stdlogicvector(X"00");
	mem(199) := To_stdlogicvector(X"00");
	mem(200) := To_stdlogicvector(X"80");
	mem(201) := To_stdlogicvector(X"C0");
	mem(202) := To_stdlogicvector(X"00");
	mem(203) := To_stdlogicvector(X"00");
	mem(204) := To_stdlogicvector(X"00");
	mem(205) := To_stdlogicvector(X"00");
	mem(206) := To_stdlogicvector(X"00");
	mem(207) := To_stdlogicvector(X"00");
	mem(208) := To_stdlogicvector(X"0A");
	mem(209) := To_stdlogicvector(X"62");
	mem(210) := To_stdlogicvector(X"00");
	mem(211) := To_stdlogicvector(X"00");
	mem(212) := To_stdlogicvector(X"00");
	mem(213) := To_stdlogicvector(X"00");
	mem(214) := To_stdlogicvector(X"00");
	mem(215) := To_stdlogicvector(X"00");
	mem(216) := To_stdlogicvector(X"0B");
	mem(217) := To_stdlogicvector(X"72");
	mem(218) := To_stdlogicvector(X"00");
	mem(219) := To_stdlogicvector(X"00");
	mem(220) := To_stdlogicvector(X"00");
	mem(221) := To_stdlogicvector(X"00");
	mem(222) := To_stdlogicvector(X"00");
	mem(223) := To_stdlogicvector(X"00");
	mem(224) := To_stdlogicvector(X"04");
	mem(225) := To_stdlogicvector(X"64");
	mem(226) := To_stdlogicvector(X"00");
	mem(227) := To_stdlogicvector(X"00");
	mem(228) := To_stdlogicvector(X"00");
	mem(229) := To_stdlogicvector(X"00");
	mem(230) := To_stdlogicvector(X"00");
	mem(231) := To_stdlogicvector(X"00");
	mem(232) := To_stdlogicvector(X"18");
	mem(233) := To_stdlogicvector(X"74");
	mem(234) := To_stdlogicvector(X"08");
	mem(235) := To_stdlogicvector(X"66");
	mem(236) := To_stdlogicvector(X"05");
	mem(237) := To_stdlogicvector(X"68");
	mem(238) := To_stdlogicvector(X"00");
	mem(239) := To_stdlogicvector(X"00");
	mem(240) := To_stdlogicvector(X"00");
	mem(241) := To_stdlogicvector(X"00");
	mem(242) := To_stdlogicvector(X"00");
	mem(243) := To_stdlogicvector(X"00");
	mem(244) := To_stdlogicvector(X"19");
	mem(245) := To_stdlogicvector(X"76");
	mem(246) := To_stdlogicvector(X"1A");
	mem(247) := To_stdlogicvector(X"78");
	mem(248) := To_stdlogicvector(X"0D");
	mem(249) := To_stdlogicvector(X"6A");
	mem(250) := To_stdlogicvector(X"00");
	mem(251) := To_stdlogicvector(X"00");
	mem(252) := To_stdlogicvector(X"00");
	mem(253) := To_stdlogicvector(X"00");
	mem(254) := To_stdlogicvector(X"00");
	mem(255) := To_stdlogicvector(X"00");
	mem(256) := To_stdlogicvector(X"1B");
	mem(257) := To_stdlogicvector(X"7A");
	mem(258) := To_stdlogicvector(X"00");
	mem(259) := To_stdlogicvector(X"00");
	mem(260) := To_stdlogicvector(X"00");
	mem(261) := To_stdlogicvector(X"00");
	mem(262) := To_stdlogicvector(X"00");
	mem(263) := To_stdlogicvector(X"00");
	mem(264) := To_stdlogicvector(X"18");
	mem(265) := To_stdlogicvector(X"6A");
	mem(266) := To_stdlogicvector(X"19");
	mem(267) := To_stdlogicvector(X"68");
	mem(268) := To_stdlogicvector(X"1A");
	mem(269) := To_stdlogicvector(X"66");
	mem(270) := To_stdlogicvector(X"1B");
	mem(271) := To_stdlogicvector(X"64");
	mem(272) := To_stdlogicvector(X"1B");
	mem(273) := To_stdlogicvector(X"7A");
	mem(274) := To_stdlogicvector(X"1B");
	mem(275) := To_stdlogicvector(X"78");
	mem(276) := To_stdlogicvector(X"1B");
	mem(277) := To_stdlogicvector(X"76");
	mem(278) := To_stdlogicvector(X"1B");
	mem(279) := To_stdlogicvector(X"74");
	mem(280) := To_stdlogicvector(X"00");
	mem(281) := To_stdlogicvector(X"00");
	mem(282) := To_stdlogicvector(X"00");
	mem(283) := To_stdlogicvector(X"00");
	mem(284) := To_stdlogicvector(X"00");
	mem(285) := To_stdlogicvector(X"00");
	mem(286) := To_stdlogicvector(X"83");
	mem(287) := To_stdlogicvector(X"14");
	mem(288) := To_stdlogicvector(X"00");
	mem(289) := To_stdlogicvector(X"00");
	mem(290) := To_stdlogicvector(X"00");
	mem(291) := To_stdlogicvector(X"00");
	mem(292) := To_stdlogicvector(X"00");
	mem(293) := To_stdlogicvector(X"00");
	mem(294) := To_stdlogicvector(X"05");
	mem(295) := To_stdlogicvector(X"17");
	mem(296) := To_stdlogicvector(X"00");
	mem(297) := To_stdlogicvector(X"00");
	mem(298) := To_stdlogicvector(X"00");
	mem(299) := To_stdlogicvector(X"00");
	mem(300) := To_stdlogicvector(X"00");
	mem(301) := To_stdlogicvector(X"00");
	mem(302) := To_stdlogicvector(X"83");
	mem(303) := To_stdlogicvector(X"14");
	mem(304) := To_stdlogicvector(X"00");
	mem(305) := To_stdlogicvector(X"00");
	mem(306) := To_stdlogicvector(X"00");
	mem(307) := To_stdlogicvector(X"00");
	mem(308) := To_stdlogicvector(X"00");
	mem(309) := To_stdlogicvector(X"00");
	mem(310) := To_stdlogicvector(X"21");
	mem(311) := To_stdlogicvector(X"16");
	mem(312) := To_stdlogicvector(X"00");
	mem(313) := To_stdlogicvector(X"00");
	mem(314) := To_stdlogicvector(X"00");
	mem(315) := To_stdlogicvector(X"00");
	mem(316) := To_stdlogicvector(X"00");
	mem(317) := To_stdlogicvector(X"00");
	mem(318) := To_stdlogicvector(X"C2");
	mem(319) := To_stdlogicvector(X"3C");
	mem(320) := To_stdlogicvector(X"01");
	mem(321) := To_stdlogicvector(X"68");
	mem(322) := To_stdlogicvector(X"04");
	mem(323) := To_stdlogicvector(X"3E");
	mem(324) := To_stdlogicvector(X"02");
	mem(325) := To_stdlogicvector(X"66");
	mem(326) := To_stdlogicvector(X"00");
	mem(327) := To_stdlogicvector(X"00");
	mem(328) := To_stdlogicvector(X"00");
	mem(329) := To_stdlogicvector(X"00");
	mem(330) := To_stdlogicvector(X"00");
	mem(331) := To_stdlogicvector(X"00");
	mem(332) := To_stdlogicvector(X"15");
	mem(333) := To_stdlogicvector(X"76");
	mem(334) := To_stdlogicvector(X"15");
	mem(335) := To_stdlogicvector(X"78");
	mem(336) := To_stdlogicvector(X"C4");
	mem(337) := To_stdlogicvector(X"16");
	mem(338) := To_stdlogicvector(X"00");
	mem(339) := To_stdlogicvector(X"68");
	mem(340) := To_stdlogicvector(X"6F");
	mem(341) := To_stdlogicvector(X"48");
	mem(342) := To_stdlogicvector(X"1E");
	mem(343) := To_stdlogicvector(X"78");
	mem(344) := To_stdlogicvector(X"72");
	mem(345) := To_stdlogicvector(X"EA");
	mem(346) := To_stdlogicvector(X"00");
	mem(347) := To_stdlogicvector(X"00");
	mem(348) := To_stdlogicvector(X"00");
	mem(349) := To_stdlogicvector(X"00");
	mem(350) := To_stdlogicvector(X"00");
	mem(351) := To_stdlogicvector(X"00");
	mem(352) := To_stdlogicvector(X"40");
	mem(353) := To_stdlogicvector(X"41");
	mem(354) := To_stdlogicvector(X"1E");
	mem(355) := To_stdlogicvector(X"7A");
	mem(356) := To_stdlogicvector(X"21");
	mem(357) := To_stdlogicvector(X"1C");
	mem(358) := To_stdlogicvector(X"00");
	mem(359) := To_stdlogicvector(X"00");
	mem(360) := To_stdlogicvector(X"00");
	mem(361) := To_stdlogicvector(X"00");
	mem(362) := To_stdlogicvector(X"00");
	mem(363) := To_stdlogicvector(X"00");
	mem(364) := To_stdlogicvector(X"9C");
	mem(365) := To_stdlogicvector(X"2D");
	mem(366) := To_stdlogicvector(X"00");
	mem(367) := To_stdlogicvector(X"00");
	mem(368) := To_stdlogicvector(X"1C");
	mem(369) := To_stdlogicvector(X"2E");
	mem(370) := To_stdlogicvector(X"00");
	mem(371) := To_stdlogicvector(X"00");
	mem(372) := To_stdlogicvector(X"16");
	mem(373) := To_stdlogicvector(X"7C");
	mem(374) := To_stdlogicvector(X"00");
	mem(375) := To_stdlogicvector(X"00");
	mem(376) := To_stdlogicvector(X"16");
	mem(377) := To_stdlogicvector(X"7E");
	mem(378) := To_stdlogicvector(X"00");
	mem(379) := To_stdlogicvector(X"00");
	mem(380) := To_stdlogicvector(X"00");
	mem(381) := To_stdlogicvector(X"00");
	mem(382) := To_stdlogicvector(X"00");
	mem(383) := To_stdlogicvector(X"00");
	mem(384) := To_stdlogicvector(X"87");
	mem(385) := To_stdlogicvector(X"1D");
	mem(386) := To_stdlogicvector(X"FD");
	mem(387) := To_stdlogicvector(X"F0");
	mem(388) := To_stdlogicvector(X"03");
	mem(389) := To_stdlogicvector(X"7C");
	mem(390) := To_stdlogicvector(X"00");
	mem(391) := To_stdlogicvector(X"62");
	mem(392) := To_stdlogicvector(X"00");
	mem(393) := To_stdlogicvector(X"64");
	mem(394) := To_stdlogicvector(X"00");
	mem(395) := To_stdlogicvector(X"66");
	mem(396) := To_stdlogicvector(X"0D");
	mem(397) := To_stdlogicvector(X"68");
	mem(398) := To_stdlogicvector(X"0D");
	mem(399) := To_stdlogicvector(X"6A");
	mem(400) := To_stdlogicvector(X"0D");
	mem(401) := To_stdlogicvector(X"6C");
	mem(402) := To_stdlogicvector(X"1C");
	mem(403) := To_stdlogicvector(X"A2");
	mem(404) := To_stdlogicvector(X"00");
	mem(405) := To_stdlogicvector(X"00");
	mem(406) := To_stdlogicvector(X"00");
	mem(407) := To_stdlogicvector(X"00");
	mem(408) := To_stdlogicvector(X"00");
	mem(409) := To_stdlogicvector(X"00");
	mem(410) := To_stdlogicvector(X"1D");
	mem(411) := To_stdlogicvector(X"B8");
	mem(412) := To_stdlogicvector(X"00");
	mem(413) := To_stdlogicvector(X"00");
	mem(414) := To_stdlogicvector(X"00");
	mem(415) := To_stdlogicvector(X"00");
	mem(416) := To_stdlogicvector(X"00");
	mem(417) := To_stdlogicvector(X"00");
	mem(418) := To_stdlogicvector(X"0C");
	mem(419) := To_stdlogicvector(X"64");
	mem(420) := To_stdlogicvector(X"0A");
	mem(421) := To_stdlogicvector(X"72");
	mem(422) := To_stdlogicvector(X"0A");
	mem(423) := To_stdlogicvector(X"74");
	mem(424) := To_stdlogicvector(X"00");
	mem(425) := To_stdlogicvector(X"00");
	mem(426) := To_stdlogicvector(X"E0");
	mem(427) := To_stdlogicvector(X"56");
	mem(428) := To_stdlogicvector(X"05");
	mem(429) := To_stdlogicvector(X"02");
	mem(430) := To_stdlogicvector(X"04");
	mem(431) := To_stdlogicvector(X"08");
	mem(432) := To_stdlogicvector(X"03");
	mem(433) := To_stdlogicvector(X"0A");
	mem(434) := To_stdlogicvector(X"03");
	mem(435) := To_stdlogicvector(X"04");
	mem(436) := To_stdlogicvector(X"01");
	mem(437) := To_stdlogicvector(X"0C");
	mem(438) := To_stdlogicvector(X"00");
	mem(439) := To_stdlogicvector(X"0E");
	mem(440) := To_stdlogicvector(X"E4");
	mem(441) := To_stdlogicvector(X"16");
	mem(442) := To_stdlogicvector(X"E6");
	mem(443) := To_stdlogicvector(X"16");
	mem(444) := To_stdlogicvector(X"20");
	mem(445) := To_stdlogicvector(X"59");
	mem(446) := To_stdlogicvector(X"01");
	mem(447) := To_stdlogicvector(X"04");
	mem(448) := To_stdlogicvector(X"E1");
	mem(449) := To_stdlogicvector(X"16");
	mem(450) := To_stdlogicvector(X"E6");
	mem(451) := To_stdlogicvector(X"16");
	mem(452) := To_stdlogicvector(X"20");
	mem(453) := To_stdlogicvector(X"59");
	mem(454) := To_stdlogicvector(X"06");
	mem(455) := To_stdlogicvector(X"0A");
	mem(456) := To_stdlogicvector(X"00");
	mem(457) := To_stdlogicvector(X"00");
	mem(458) := To_stdlogicvector(X"00");
	mem(459) := To_stdlogicvector(X"00");
	mem(460) := To_stdlogicvector(X"00");
	mem(461) := To_stdlogicvector(X"00");
	mem(462) := To_stdlogicvector(X"2A");
	mem(463) := To_stdlogicvector(X"19");
	mem(464) := To_stdlogicvector(X"00");
	mem(465) := To_stdlogicvector(X"00");
	mem(466) := To_stdlogicvector(X"02");
	mem(467) := To_stdlogicvector(X"02");
	mem(468) := To_stdlogicvector(X"E6");
	mem(469) := To_stdlogicvector(X"16");
	mem(470) := To_stdlogicvector(X"04");
	mem(471) := To_stdlogicvector(X"0E");
	mem(472) := To_stdlogicvector(X"E3");
	mem(473) := To_stdlogicvector(X"16");
	mem(474) := To_stdlogicvector(X"00");
	mem(475) := To_stdlogicvector(X"00");
	mem(476) := To_stdlogicvector(X"00");
	mem(477) := To_stdlogicvector(X"00");
	mem(478) := To_stdlogicvector(X"00");
	mem(479) := To_stdlogicvector(X"00");
	mem(480) := To_stdlogicvector(X"C4");
	mem(481) := To_stdlogicvector(X"16");
	mem(482) := To_stdlogicvector(X"00");
	mem(483) := To_stdlogicvector(X"00");
	mem(484) := To_stdlogicvector(X"00");
	mem(485) := To_stdlogicvector(X"00");
	mem(486) := To_stdlogicvector(X"00");
	mem(487) := To_stdlogicvector(X"00");
	mem(488) := To_stdlogicvector(X"0A");
	mem(489) := To_stdlogicvector(X"76");
	mem(490) := To_stdlogicvector(X"18");
	mem(491) := To_stdlogicvector(X"72");
	mem(492) := To_stdlogicvector(X"19");
	mem(493) := To_stdlogicvector(X"74");
	mem(494) := To_stdlogicvector(X"1A");
	mem(495) := To_stdlogicvector(X"76");
	mem(496) := To_stdlogicvector(X"2F");
	mem(497) := To_stdlogicvector(X"E2");
	mem(498) := To_stdlogicvector(X"40");
	mem(499) := To_stdlogicvector(X"C0");
	mem(500) := To_stdlogicvector(X"00");
	mem(501) := To_stdlogicvector(X"00");
	mem(502) := To_stdlogicvector(X"0F");
	mem(503) := To_stdlogicvector(X"70");
	mem(504) := To_stdlogicvector(X"AD");
	mem(505) := To_stdlogicvector(X"BE");
	mem(506) := To_stdlogicvector(X"42");
	mem(507) := To_stdlogicvector(X"02");
	mem(508) := To_stdlogicvector(X"EB");
	mem(509) := To_stdlogicvector(X"DE");
	mem(510) := To_stdlogicvector(X"AF");
	mem(511) := To_stdlogicvector(X"1E");
	mem(512) := To_stdlogicvector(X"2D");
	mem(513) := To_stdlogicvector(X"D2");
	mem(514) := To_stdlogicvector(X"42");
	mem(515) := To_stdlogicvector(X"00");
	mem(516) := To_stdlogicvector(X"ED");
	mem(517) := To_stdlogicvector(X"F0");
	mem(518) := To_stdlogicvector(X"06");
	mem(519) := To_stdlogicvector(X"B0");
	mem(520) := To_stdlogicvector(X"0F");
	mem(521) := To_stdlogicvector(X"60");
	mem(522) := To_stdlogicvector(X"DD");
	mem(523) := To_stdlogicvector(X"DD");
	mem(524) := To_stdlogicvector(X"00");
	mem(525) := To_stdlogicvector(X"00");
	mem(526) := To_stdlogicvector(X"0D");
	mem(527) := To_stdlogicvector(X"60");
	mem(528) := To_stdlogicvector(X"CA");
	mem(529) := To_stdlogicvector(X"D0");
	mem(530) := To_stdlogicvector(X"0B");
	mem(531) := To_stdlogicvector(X"F0");
	mem(532) := To_stdlogicvector(X"FF");
	mem(533) := To_stdlogicvector(X"FF");
	mem(534) := To_stdlogicvector(X"10");
	mem(535) := To_stdlogicvector(X"10");
	mem(536) := To_stdlogicvector(X"34");
	mem(537) := To_stdlogicvector(X"12");
	mem(538) := To_stdlogicvector(X"21");
	mem(539) := To_stdlogicvector(X"89");
	mem(540) := To_stdlogicvector(X"99");
	mem(541) := To_stdlogicvector(X"99");
	mem(542) := To_stdlogicvector(X"CC");
	mem(543) := To_stdlogicvector(X"CC");
	mem(544) := To_stdlogicvector(X"69");
	mem(545) := To_stdlogicvector(X"69");
	mem(546) := To_stdlogicvector(X"11");
	mem(547) := To_stdlogicvector(X"BA");
	mem(548) := To_stdlogicvector(X"88");
	mem(549) := To_stdlogicvector(X"88");
	mem(550) := To_stdlogicvector(X"CD");
	mem(551) := To_stdlogicvector(X"AB");
	mem(552) := To_stdlogicvector(X"10");
	mem(553) := To_stdlogicvector(X"01");
	mem(554) := To_stdlogicvector(X"BA");
	mem(555) := To_stdlogicvector(X"AB");
	mem(556) := To_stdlogicvector(X"22");
	mem(557) := To_stdlogicvector(X"02");
	mem(558) := To_stdlogicvector(X"0C");
	mem(559) := To_stdlogicvector(X"02");
	mem(560) := To_stdlogicvector(X"00");
	mem(561) := To_stdlogicvector(X"00");
	mem(562) := To_stdlogicvector(X"50");
	mem(563) := To_stdlogicvector(X"02");
	mem(564) := To_stdlogicvector(X"00");
	mem(565) := To_stdlogicvector(X"00");
	mem(566) := To_stdlogicvector(X"00");
	mem(567) := To_stdlogicvector(X"00");
	mem(568) := To_stdlogicvector(X"00");
	mem(569) := To_stdlogicvector(X"00");
	mem(570) := To_stdlogicvector(X"2E");
	mem(571) := To_stdlogicvector(X"19");
	mem(572) := To_stdlogicvector(X"C0");
	mem(573) := To_stdlogicvector(X"C1");
	mem(574) := To_stdlogicvector(X"07");
	mem(575) := To_stdlogicvector(X"6A");
	mem(576) := To_stdlogicvector(X"C0");
	mem(577) := To_stdlogicvector(X"C1");
	mem(578) := To_stdlogicvector(X"0D");
	mem(579) := To_stdlogicvector(X"62");
	mem(580) := To_stdlogicvector(X"0D");
	mem(581) := To_stdlogicvector(X"64");
	mem(582) := To_stdlogicvector(X"0D");
	mem(583) := To_stdlogicvector(X"66");
	mem(584) := To_stdlogicvector(X"0D");
	mem(585) := To_stdlogicvector(X"68");
	mem(586) := To_stdlogicvector(X"0D");
	mem(587) := To_stdlogicvector(X"6A");
	mem(588) := To_stdlogicvector(X"0D");
	mem(589) := To_stdlogicvector(X"6C");
	mem(590) := To_stdlogicvector(X"C0");
	mem(591) := To_stdlogicvector(X"C1");
	mem(592) := To_stdlogicvector(X"6B");
	mem(593) := To_stdlogicvector(X"E0");
	mem(594) := To_stdlogicvector(X"60");
	mem(595) := To_stdlogicvector(X"52");
	mem(596) := To_stdlogicvector(X"A0");
	mem(597) := To_stdlogicvector(X"54");
	mem(598) := To_stdlogicvector(X"E0");
	mem(599) := To_stdlogicvector(X"56");
	mem(600) := To_stdlogicvector(X"ED");
	mem(601) := To_stdlogicvector(X"16");
	mem(602) := To_stdlogicvector(X"AB");
	mem(603) := To_stdlogicvector(X"14");
	mem(604) := To_stdlogicvector(X"83");
	mem(605) := To_stdlogicvector(X"12");
	mem(606) := To_stdlogicvector(X"63");
	mem(607) := To_stdlogicvector(X"18");
	mem(608) := To_stdlogicvector(X"A3");
	mem(609) := To_stdlogicvector(X"D4");
	mem(610) := To_stdlogicvector(X"FF");
	mem(611) := To_stdlogicvector(X"9A");
	mem(612) := To_stdlogicvector(X"AF");
	mem(613) := To_stdlogicvector(X"56");
	mem(614) := To_stdlogicvector(X"00");
	mem(615) := To_stdlogicvector(X"00");
	mem(616) := To_stdlogicvector(X"00");
	mem(617) := To_stdlogicvector(X"00");
	mem(618) := To_stdlogicvector(X"C3");
	mem(619) := To_stdlogicvector(X"1A");
	mem(620) := To_stdlogicvector(X"25");
	mem(621) := To_stdlogicvector(X"13");
	mem(622) := To_stdlogicvector(X"2A");
	mem(623) := To_stdlogicvector(X"13");
	mem(624) := To_stdlogicvector(X"2E");
	mem(625) := To_stdlogicvector(X"13");
	mem(626) := To_stdlogicvector(X"7F");
	mem(627) := To_stdlogicvector(X"54");
	mem(628) := To_stdlogicvector(X"00");
	mem(629) := To_stdlogicvector(X"74");
	mem(630) := To_stdlogicvector(X"00");
	mem(631) := To_stdlogicvector(X"7A");
	mem(632) := To_stdlogicvector(X"22");
	mem(633) := To_stdlogicvector(X"10");
	mem(634) := To_stdlogicvector(X"00");
	mem(635) := To_stdlogicvector(X"74");
	mem(636) := To_stdlogicvector(X"3E");
	mem(637) := To_stdlogicvector(X"10");
	mem(638) := To_stdlogicvector(X"03");
	mem(639) := To_stdlogicvector(X"66");
	mem(640) := To_stdlogicvector(X"02");
	mem(641) := To_stdlogicvector(X"66");
	mem(642) := To_stdlogicvector(X"03");
	mem(643) := To_stdlogicvector(X"76");
	mem(644) := To_stdlogicvector(X"04");
	mem(645) := To_stdlogicvector(X"66");
	mem(646) := To_stdlogicvector(X"EB");
	mem(647) := To_stdlogicvector(X"18");
	mem(648) := To_stdlogicvector(X"05");
	mem(649) := To_stdlogicvector(X"66");
	mem(650) := To_stdlogicvector(X"11");
	mem(651) := To_stdlogicvector(X"D9");
	mem(652) := To_stdlogicvector(X"E7");
	mem(653) := To_stdlogicvector(X"1A");
	mem(654) := To_stdlogicvector(X"06");
	mem(655) := To_stdlogicvector(X"A2");
	mem(656) := To_stdlogicvector(X"6C");
	mem(657) := To_stdlogicvector(X"1B");
	mem(658) := To_stdlogicvector(X"2C");
	mem(659) := To_stdlogicvector(X"13");
	mem(660) := To_stdlogicvector(X"EC");
	mem(661) := To_stdlogicvector(X"14");
	mem(662) := To_stdlogicvector(X"07");
	mem(663) := To_stdlogicvector(X"72");
	mem(664) := To_stdlogicvector(X"07");
	mem(665) := To_stdlogicvector(X"74");
	mem(666) := To_stdlogicvector(X"07");
	mem(667) := To_stdlogicvector(X"76");
	mem(668) := To_stdlogicvector(X"07");
	mem(669) := To_stdlogicvector(X"78");
	mem(670) := To_stdlogicvector(X"07");
	mem(671) := To_stdlogicvector(X"7A");
	mem(672) := To_stdlogicvector(X"60");
	mem(673) := To_stdlogicvector(X"1A");
	mem(674) := To_stdlogicvector(X"E0");
	mem(675) := To_stdlogicvector(X"1C");
	mem(676) := To_stdlogicvector(X"20");
	mem(677) := To_stdlogicvector(X"1F");
	mem(678) := To_stdlogicvector(X"60");
	mem(679) := To_stdlogicvector(X"52");
	mem(680) := To_stdlogicvector(X"E0");
	mem(681) := To_stdlogicvector(X"56");
	mem(682) := To_stdlogicvector(X"20");
	mem(683) := To_stdlogicvector(X"59");
	mem(684) := To_stdlogicvector(X"68");
	mem(685) := To_stdlogicvector(X"12");
	mem(686) := To_stdlogicvector(X"E2");
	mem(687) := To_stdlogicvector(X"16");
	mem(688) := To_stdlogicvector(X"22");
	mem(689) := To_stdlogicvector(X"19");
	mem(690) := To_stdlogicvector(X"01");
	mem(691) := To_stdlogicvector(X"02");
	mem(692) := To_stdlogicvector(X"E1");
	mem(693) := To_stdlogicvector(X"16");
	mem(694) := To_stdlogicvector(X"69");
	mem(695) := To_stdlogicvector(X"12");
	mem(696) := To_stdlogicvector(X"0C");
	mem(697) := To_stdlogicvector(X"08");
	mem(698) := To_stdlogicvector(X"21");
	mem(699) := To_stdlogicvector(X"19");
	mem(700) := To_stdlogicvector(X"07");
	mem(701) := To_stdlogicvector(X"60");
	mem(702) := To_stdlogicvector(X"9A");
	mem(703) := To_stdlogicvector(X"E1");
	mem(704) := To_stdlogicvector(X"18");
	mem(705) := To_stdlogicvector(X"64");
	mem(706) := To_stdlogicvector(X"19");
	mem(707) := To_stdlogicvector(X"6C");
	mem(708) := To_stdlogicvector(X"1A");
	mem(709) := To_stdlogicvector(X"6E");
	mem(710) := To_stdlogicvector(X"30");
	mem(711) := To_stdlogicvector(X"E0");
	mem(712) := To_stdlogicvector(X"E0");
	mem(713) := To_stdlogicvector(X"56");
	mem(714) := To_stdlogicvector(X"20");
	mem(715) := To_stdlogicvector(X"59");
	mem(716) := To_stdlogicvector(X"00");
	mem(717) := To_stdlogicvector(X"00");
	mem(718) := To_stdlogicvector(X"E2");
	mem(719) := To_stdlogicvector(X"16");
	mem(720) := To_stdlogicvector(X"23");
	mem(721) := To_stdlogicvector(X"19");
	mem(722) := To_stdlogicvector(X"08");
	mem(723) := To_stdlogicvector(X"62");
	mem(724) := To_stdlogicvector(X"01");
	mem(725) := To_stdlogicvector(X"08");
	mem(726) := To_stdlogicvector(X"E1");
	mem(727) := To_stdlogicvector(X"16");
	mem(728) := To_stdlogicvector(X"09");
	mem(729) := To_stdlogicvector(X"62");
	mem(730) := To_stdlogicvector(X"01");
	mem(731) := To_stdlogicvector(X"04");
	mem(732) := To_stdlogicvector(X"21");
	mem(733) := To_stdlogicvector(X"19");
	mem(734) := To_stdlogicvector(X"0A");
	mem(735) := To_stdlogicvector(X"A2");
	mem(736) := To_stdlogicvector(X"01");
	mem(737) := To_stdlogicvector(X"0C");
	mem(738) := To_stdlogicvector(X"E1");
	mem(739) := To_stdlogicvector(X"16");
	mem(740) := To_stdlogicvector(X"06");
	mem(741) := To_stdlogicvector(X"A2");
	mem(742) := To_stdlogicvector(X"01");
	mem(743) := To_stdlogicvector(X"0C");
	mem(744) := To_stdlogicvector(X"21");
	mem(745) := To_stdlogicvector(X"19");
	mem(746) := To_stdlogicvector(X"20");
	mem(747) := To_stdlogicvector(X"52");
	mem(748) := To_stdlogicvector(X"1D");
	mem(749) := To_stdlogicvector(X"E2");
	mem(750) := To_stdlogicvector(X"01");
	mem(751) := To_stdlogicvector(X"02");
	mem(752) := To_stdlogicvector(X"E1");
	mem(753) := To_stdlogicvector(X"16");
	mem(754) := To_stdlogicvector(X"0B");
	mem(755) := To_stdlogicvector(X"76");
	mem(756) := To_stdlogicvector(X"0C");
	mem(757) := To_stdlogicvector(X"78");
	mem(758) := To_stdlogicvector(X"60");
	mem(759) := To_stdlogicvector(X"52");
	mem(760) := To_stdlogicvector(X"60");
	mem(761) := To_stdlogicvector(X"5B");
	mem(762) := To_stdlogicvector(X"7F");
	mem(763) := To_stdlogicvector(X"12");
	mem(764) := To_stdlogicvector(X"02");
	mem(765) := To_stdlogicvector(X"08");
	mem(766) := To_stdlogicvector(X"61");
	mem(767) := To_stdlogicvector(X"1B");
	mem(768) := To_stdlogicvector(X"79");
	mem(769) := To_stdlogicvector(X"12");
	mem(770) := To_stdlogicvector(X"45");
	mem(771) := To_stdlogicvector(X"1A");
	mem(772) := To_stdlogicvector(X"00");
	mem(773) := To_stdlogicvector(X"00");
	mem(774) := To_stdlogicvector(X"00");
	mem(775) := To_stdlogicvector(X"00");
	mem(776) := To_stdlogicvector(X"00");
	mem(777) := To_stdlogicvector(X"00");
	mem(778) := To_stdlogicvector(X"0D");
	mem(779) := To_stdlogicvector(X"7A");
	mem(780) := To_stdlogicvector(X"60");
	mem(781) := To_stdlogicvector(X"11");
	mem(782) := To_stdlogicvector(X"60");
	mem(783) := To_stdlogicvector(X"5B");
	mem(784) := To_stdlogicvector(X"02");
	mem(785) := To_stdlogicvector(X"E2");
	mem(786) := To_stdlogicvector(X"40");
	mem(787) := To_stdlogicvector(X"C0");
	mem(788) := To_stdlogicvector(X"61");
	mem(789) := To_stdlogicvector(X"1B");
	mem(790) := To_stdlogicvector(X"05");
	mem(791) := To_stdlogicvector(X"1A");
	mem(792) := To_stdlogicvector(X"6D");
	mem(793) := To_stdlogicvector(X"E1");
	mem(794) := To_stdlogicvector(X"00");
	mem(795) := To_stdlogicvector(X"00");
	mem(796) := To_stdlogicvector(X"00");
	mem(797) := To_stdlogicvector(X"00");
	mem(798) := To_stdlogicvector(X"00");
	mem(799) := To_stdlogicvector(X"00");
	mem(800) := To_stdlogicvector(X"03");
	mem(801) := To_stdlogicvector(X"62");
	mem(802) := To_stdlogicvector(X"02");
	mem(803) := To_stdlogicvector(X"E0");
	mem(804) := To_stdlogicvector(X"00");
	mem(805) := To_stdlogicvector(X"7A");
	mem(806) := To_stdlogicvector(X"10");
	mem(807) := To_stdlogicvector(X"0E");
	mem(808) := To_stdlogicvector(X"00");
	mem(809) := To_stdlogicvector(X"00");
	mem(810) := To_stdlogicvector(X"00");
	mem(811) := To_stdlogicvector(X"00");
	mem(812) := To_stdlogicvector(X"DA");
	mem(813) := To_stdlogicvector(X"AB");
	mem(814) := To_stdlogicvector(X"00");
	mem(815) := To_stdlogicvector(X"00");
	mem(816) := To_stdlogicvector(X"4D");
	mem(817) := To_stdlogicvector(X"9A");
	mem(818) := To_stdlogicvector(X"AC");
	mem(819) := To_stdlogicvector(X"3D");
	mem(820) := To_stdlogicvector(X"44");
	mem(821) := To_stdlogicvector(X"03");
	mem(822) := To_stdlogicvector(X"DD");
	mem(823) := To_stdlogicvector(X"FA");
	mem(824) := To_stdlogicvector(X"03");
	mem(825) := To_stdlogicvector(X"FB");
	mem(826) := To_stdlogicvector(X"11");
	mem(827) := To_stdlogicvector(X"01");
	mem(828) := To_stdlogicvector(X"38");
	mem(829) := To_stdlogicvector(X"03");
	mem(830) := To_stdlogicvector(X"0F");
	mem(831) := To_stdlogicvector(X"F0");
	mem(832) := To_stdlogicvector(X"0F");
	mem(833) := To_stdlogicvector(X"F0");
	mem(834) := To_stdlogicvector(X"EE");
	mem(835) := To_stdlogicvector(X"0F");
	mem(836) := To_stdlogicvector(X"6C");
	mem(837) := To_stdlogicvector(X"27");
	mem(838) := To_stdlogicvector(X"48");
	mem(839) := To_stdlogicvector(X"03");
	mem(840) := To_stdlogicvector(X"E0");
	mem(841) := To_stdlogicvector(X"5F");
	mem(842) := To_stdlogicvector(X"A0");
	mem(843) := To_stdlogicvector(X"5D");
	mem(844) := To_stdlogicvector(X"60");
	mem(845) := To_stdlogicvector(X"5B");
	mem(846) := To_stdlogicvector(X"20");
	mem(847) := To_stdlogicvector(X"59");
	mem(848) := To_stdlogicvector(X"E0");
	mem(849) := To_stdlogicvector(X"56");
	mem(850) := To_stdlogicvector(X"A0");
	mem(851) := To_stdlogicvector(X"54");
	mem(852) := To_stdlogicvector(X"60");
	mem(853) := To_stdlogicvector(X"52");
	mem(854) := To_stdlogicvector(X"20");
	mem(855) := To_stdlogicvector(X"50");
	mem(856) := To_stdlogicvector(X"B6");
	mem(857) := To_stdlogicvector(X"E0");
	mem(858) := To_stdlogicvector(X"C4");
	mem(859) := To_stdlogicvector(X"E2");
	mem(860) := To_stdlogicvector(X"0B");
	mem(861) := To_stdlogicvector(X"64");
	mem(862) := To_stdlogicvector(X"08");
	mem(863) := To_stdlogicvector(X"66");
	mem(864) := To_stdlogicvector(X"40");
	mem(865) := To_stdlogicvector(X"74");
	mem(866) := To_stdlogicvector(X"B9");
	mem(867) := To_stdlogicvector(X"14");
	mem(868) := To_stdlogicvector(X"62");
	mem(869) := To_stdlogicvector(X"12");
	mem(870) := To_stdlogicvector(X"FF");
	mem(871) := To_stdlogicvector(X"16");
	mem(872) := To_stdlogicvector(X"FB");
	mem(873) := To_stdlogicvector(X"03");
	mem(874) := To_stdlogicvector(X"BC");
	mem(875) := To_stdlogicvector(X"E8");
	mem(876) := To_stdlogicvector(X"08");
	mem(877) := To_stdlogicvector(X"64");
	mem(878) := To_stdlogicvector(X"84");
	mem(879) := To_stdlogicvector(X"18");
	mem(880) := To_stdlogicvector(X"0B");
	mem(881) := To_stdlogicvector(X"66");
	mem(882) := To_stdlogicvector(X"60");
	mem(883) := To_stdlogicvector(X"52");
	mem(884) := To_stdlogicvector(X"A0");
	mem(885) := To_stdlogicvector(X"54");
	mem(886) := To_stdlogicvector(X"7D");
	mem(887) := To_stdlogicvector(X"48");
	mem(888) := To_stdlogicvector(X"44");
	mem(889) := To_stdlogicvector(X"1D");
	mem(890) := To_stdlogicvector(X"80");
	mem(891) := To_stdlogicvector(X"77");
	mem(892) := To_stdlogicvector(X"FE");
	mem(893) := To_stdlogicvector(X"16");
	mem(894) := To_stdlogicvector(X"55");
	mem(895) := To_stdlogicvector(X"48");
	mem(896) := To_stdlogicvector(X"60");
	mem(897) := To_stdlogicvector(X"1A");
	mem(898) := To_stdlogicvector(X"F9");
	mem(899) := To_stdlogicvector(X"07");
	mem(900) := To_stdlogicvector(X"AF");
	mem(901) := To_stdlogicvector(X"E8");
	mem(902) := To_stdlogicvector(X"08");
	mem(903) := To_stdlogicvector(X"64");
	mem(904) := To_stdlogicvector(X"84");
	mem(905) := To_stdlogicvector(X"18");
	mem(906) := To_stdlogicvector(X"84");
	mem(907) := To_stdlogicvector(X"18");
	mem(908) := To_stdlogicvector(X"0B");
	mem(909) := To_stdlogicvector(X"66");
	mem(910) := To_stdlogicvector(X"60");
	mem(911) := To_stdlogicvector(X"52");
	mem(912) := To_stdlogicvector(X"A0");
	mem(913) := To_stdlogicvector(X"54");
	mem(914) := To_stdlogicvector(X"6F");
	mem(915) := To_stdlogicvector(X"48");
	mem(916) := To_stdlogicvector(X"44");
	mem(917) := To_stdlogicvector(X"1D");
	mem(918) := To_stdlogicvector(X"80");
	mem(919) := To_stdlogicvector(X"77");
	mem(920) := To_stdlogicvector(X"FB");
	mem(921) := To_stdlogicvector(X"16");
	mem(922) := To_stdlogicvector(X"53");
	mem(923) := To_stdlogicvector(X"48");
	mem(924) := To_stdlogicvector(X"60");
	mem(925) := To_stdlogicvector(X"1A");
	mem(926) := To_stdlogicvector(X"F9");
	mem(927) := To_stdlogicvector(X"07");
	mem(928) := To_stdlogicvector(X"A1");
	mem(929) := To_stdlogicvector(X"E6");
	mem(930) := To_stdlogicvector(X"08");
	mem(931) := To_stdlogicvector(X"68");
	mem(932) := To_stdlogicvector(X"C4");
	mem(933) := To_stdlogicvector(X"18");
	mem(934) := To_stdlogicvector(X"A0");
	mem(935) := To_stdlogicvector(X"5D");
	mem(936) := To_stdlogicvector(X"02");
	mem(937) := To_stdlogicvector(X"62");
	mem(938) := To_stdlogicvector(X"03");
	mem(939) := To_stdlogicvector(X"64");
	mem(940) := To_stdlogicvector(X"62");
	mem(941) := To_stdlogicvector(X"48");
	mem(942) := To_stdlogicvector(X"44");
	mem(943) := To_stdlogicvector(X"1F");
	mem(944) := To_stdlogicvector(X"C0");
	mem(945) := To_stdlogicvector(X"6D");
	mem(946) := To_stdlogicvector(X"47");
	mem(947) := To_stdlogicvector(X"48");
	mem(948) := To_stdlogicvector(X"02");
	mem(949) := To_stdlogicvector(X"72");
	mem(950) := To_stdlogicvector(X"03");
	mem(951) := To_stdlogicvector(X"74");
	mem(952) := To_stdlogicvector(X"00");
	mem(953) := To_stdlogicvector(X"62");
	mem(954) := To_stdlogicvector(X"01");
	mem(955) := To_stdlogicvector(X"64");
	mem(956) := To_stdlogicvector(X"5A");
	mem(957) := To_stdlogicvector(X"48");
	mem(958) := To_stdlogicvector(X"43");
	mem(959) := To_stdlogicvector(X"1B");
	mem(960) := To_stdlogicvector(X"40");
	mem(961) := To_stdlogicvector(X"6F");
	mem(962) := To_stdlogicvector(X"87");
	mem(963) := To_stdlogicvector(X"1D");
	mem(964) := To_stdlogicvector(X"40");
	mem(965) := To_stdlogicvector(X"7D");
	mem(966) := To_stdlogicvector(X"31");
	mem(967) := To_stdlogicvector(X"48");
	mem(968) := To_stdlogicvector(X"60");
	mem(969) := To_stdlogicvector(X"1E");
	mem(970) := To_stdlogicvector(X"03");
	mem(971) := To_stdlogicvector(X"08");
	mem(972) := To_stdlogicvector(X"00");
	mem(973) := To_stdlogicvector(X"72");
	mem(974) := To_stdlogicvector(X"01");
	mem(975) := To_stdlogicvector(X"74");
	mem(976) := To_stdlogicvector(X"EB");
	mem(977) := To_stdlogicvector(X"0F");
	mem(978) := To_stdlogicvector(X"60");
	mem(979) := To_stdlogicvector(X"52");
	mem(980) := To_stdlogicvector(X"00");
	mem(981) := To_stdlogicvector(X"72");
	mem(982) := To_stdlogicvector(X"02");
	mem(983) := To_stdlogicvector(X"72");
	mem(984) := To_stdlogicvector(X"01");
	mem(985) := To_stdlogicvector(X"72");
	mem(986) := To_stdlogicvector(X"03");
	mem(987) := To_stdlogicvector(X"72");
	mem(988) := To_stdlogicvector(X"83");
	mem(989) := To_stdlogicvector(X"E6");
	mem(990) := To_stdlogicvector(X"08");
	mem(991) := To_stdlogicvector(X"68");
	mem(992) := To_stdlogicvector(X"04");
	mem(993) := To_stdlogicvector(X"19");
	mem(994) := To_stdlogicvector(X"C4");
	mem(995) := To_stdlogicvector(X"18");
	mem(996) := To_stdlogicvector(X"A0");
	mem(997) := To_stdlogicvector(X"5D");
	mem(998) := To_stdlogicvector(X"02");
	mem(999) := To_stdlogicvector(X"62");
	mem(1000) := To_stdlogicvector(X"03");
	mem(1001) := To_stdlogicvector(X"64");
	mem(1002) := To_stdlogicvector(X"43");
	mem(1003) := To_stdlogicvector(X"48");
	mem(1004) := To_stdlogicvector(X"43");
	mem(1005) := To_stdlogicvector(X"1F");
	mem(1006) := To_stdlogicvector(X"C0");
	mem(1007) := To_stdlogicvector(X"6D");
	mem(1008) := To_stdlogicvector(X"10");
	mem(1009) := To_stdlogicvector(X"48");
	mem(1010) := To_stdlogicvector(X"02");
	mem(1011) := To_stdlogicvector(X"72");
	mem(1012) := To_stdlogicvector(X"03");
	mem(1013) := To_stdlogicvector(X"74");
	mem(1014) := To_stdlogicvector(X"00");
	mem(1015) := To_stdlogicvector(X"62");
	mem(1016) := To_stdlogicvector(X"01");
	mem(1017) := To_stdlogicvector(X"64");
	mem(1018) := To_stdlogicvector(X"3B");
	mem(1019) := To_stdlogicvector(X"48");
	mem(1020) := To_stdlogicvector(X"44");
	mem(1021) := To_stdlogicvector(X"1B");
	mem(1022) := To_stdlogicvector(X"40");
	mem(1023) := To_stdlogicvector(X"6F");
	mem(1024) := To_stdlogicvector(X"87");
	mem(1025) := To_stdlogicvector(X"1D");
	mem(1026) := To_stdlogicvector(X"40");
	mem(1027) := To_stdlogicvector(X"7D");
	mem(1028) := To_stdlogicvector(X"1E");
	mem(1029) := To_stdlogicvector(X"48");
	mem(1030) := To_stdlogicvector(X"60");
	mem(1031) := To_stdlogicvector(X"1E");
	mem(1032) := To_stdlogicvector(X"03");
	mem(1033) := To_stdlogicvector(X"08");
	mem(1034) := To_stdlogicvector(X"00");
	mem(1035) := To_stdlogicvector(X"72");
	mem(1036) := To_stdlogicvector(X"01");
	mem(1037) := To_stdlogicvector(X"74");
	mem(1038) := To_stdlogicvector(X"EB");
	mem(1039) := To_stdlogicvector(X"0F");
	mem(1040) := To_stdlogicvector(X"34");
	mem(1041) := To_stdlogicvector(X"0E");
	mem(1042) := To_stdlogicvector(X"71");
	mem(1043) := To_stdlogicvector(X"1A");
	mem(1044) := To_stdlogicvector(X"02");
	mem(1045) := To_stdlogicvector(X"04");
	mem(1046) := To_stdlogicvector(X"61");
	mem(1047) := To_stdlogicvector(X"12");
	mem(1048) := To_stdlogicvector(X"07");
	mem(1049) := To_stdlogicvector(X"0E");
	mem(1050) := To_stdlogicvector(X"B1");
	mem(1051) := To_stdlogicvector(X"1A");
	mem(1052) := To_stdlogicvector(X"03");
	mem(1053) := To_stdlogicvector(X"04");
	mem(1054) := To_stdlogicvector(X"A1");
	mem(1055) := To_stdlogicvector(X"14");
	mem(1056) := To_stdlogicvector(X"60");
	mem(1057) := To_stdlogicvector(X"52");
	mem(1058) := To_stdlogicvector(X"02");
	mem(1059) := To_stdlogicvector(X"0E");
	mem(1060) := To_stdlogicvector(X"60");
	mem(1061) := To_stdlogicvector(X"52");
	mem(1062) := To_stdlogicvector(X"7F");
	mem(1063) := To_stdlogicvector(X"12");
	mem(1064) := To_stdlogicvector(X"C0");
	mem(1065) := To_stdlogicvector(X"C1");
	mem(1066) := To_stdlogicvector(X"B1");
	mem(1067) := To_stdlogicvector(X"1A");
	mem(1068) := To_stdlogicvector(X"02");
	mem(1069) := To_stdlogicvector(X"04");
	mem(1070) := To_stdlogicvector(X"A1");
	mem(1071) := To_stdlogicvector(X"14");
	mem(1072) := To_stdlogicvector(X"07");
	mem(1073) := To_stdlogicvector(X"0E");
	mem(1074) := To_stdlogicvector(X"71");
	mem(1075) := To_stdlogicvector(X"1A");
	mem(1076) := To_stdlogicvector(X"03");
	mem(1077) := To_stdlogicvector(X"04");
	mem(1078) := To_stdlogicvector(X"61");
	mem(1079) := To_stdlogicvector(X"12");
	mem(1080) := To_stdlogicvector(X"A0");
	mem(1081) := To_stdlogicvector(X"54");
	mem(1082) := To_stdlogicvector(X"02");
	mem(1083) := To_stdlogicvector(X"0E");
	mem(1084) := To_stdlogicvector(X"60");
	mem(1085) := To_stdlogicvector(X"52");
	mem(1086) := To_stdlogicvector(X"7F");
	mem(1087) := To_stdlogicvector(X"12");
	mem(1088) := To_stdlogicvector(X"C0");
	mem(1089) := To_stdlogicvector(X"C1");
	mem(1090) := To_stdlogicvector(X"06");
	mem(1091) := To_stdlogicvector(X"76");
	mem(1092) := To_stdlogicvector(X"71");
	mem(1093) := To_stdlogicvector(X"16");
	mem(1094) := To_stdlogicvector(X"0B");
	mem(1095) := To_stdlogicvector(X"04");
	mem(1096) := To_stdlogicvector(X"A0");
	mem(1097) := To_stdlogicvector(X"16");
	mem(1098) := To_stdlogicvector(X"06");
	mem(1099) := To_stdlogicvector(X"04");
	mem(1100) := To_stdlogicvector(X"0D");
	mem(1101) := To_stdlogicvector(X"66");
	mem(1102) := To_stdlogicvector(X"71");
	mem(1103) := To_stdlogicvector(X"16");
	mem(1104) := To_stdlogicvector(X"06");
	mem(1105) := To_stdlogicvector(X"04");
	mem(1106) := To_stdlogicvector(X"61");
	mem(1107) := To_stdlogicvector(X"12");
	mem(1108) := To_stdlogicvector(X"BF");
	mem(1109) := To_stdlogicvector(X"14");
	mem(1110) := To_stdlogicvector(X"0B");
	mem(1111) := To_stdlogicvector(X"0E");
	mem(1112) := To_stdlogicvector(X"61");
	mem(1113) := To_stdlogicvector(X"14");
	mem(1114) := To_stdlogicvector(X"60");
	mem(1115) := To_stdlogicvector(X"52");
	mem(1116) := To_stdlogicvector(X"08");
	mem(1117) := To_stdlogicvector(X"0E");
	mem(1118) := To_stdlogicvector(X"B1");
	mem(1119) := To_stdlogicvector(X"16");
	mem(1120) := To_stdlogicvector(X"04");
	mem(1121) := To_stdlogicvector(X"04");
	mem(1122) := To_stdlogicvector(X"A1");
	mem(1123) := To_stdlogicvector(X"12");
	mem(1124) := To_stdlogicvector(X"A0");
	mem(1125) := To_stdlogicvector(X"54");
	mem(1126) := To_stdlogicvector(X"AF");
	mem(1127) := To_stdlogicvector(X"14");
	mem(1128) := To_stdlogicvector(X"02");
	mem(1129) := To_stdlogicvector(X"0E");
	mem(1130) := To_stdlogicvector(X"60");
	mem(1131) := To_stdlogicvector(X"52");
	mem(1132) := To_stdlogicvector(X"7F");
	mem(1133) := To_stdlogicvector(X"12");
	mem(1134) := To_stdlogicvector(X"06");
	mem(1135) := To_stdlogicvector(X"66");
	mem(1136) := To_stdlogicvector(X"C0");
	mem(1137) := To_stdlogicvector(X"C1");
	mem(1138) := To_stdlogicvector(X"A4");
	mem(1139) := To_stdlogicvector(X"DA");
	mem(1140) := To_stdlogicvector(X"45");
	mem(1141) := To_stdlogicvector(X"1A");
	mem(1142) := To_stdlogicvector(X"61");
	mem(1143) := To_stdlogicvector(X"DB");
	mem(1144) := To_stdlogicvector(X"C0");
	mem(1145) := To_stdlogicvector(X"C1");
	mem(1146) := To_stdlogicvector(X"34");
	mem(1147) := To_stdlogicvector(X"E2");
	mem(1148) := To_stdlogicvector(X"08");
	mem(1149) := To_stdlogicvector(X"68");
	mem(1150) := To_stdlogicvector(X"04");
	mem(1151) := To_stdlogicvector(X"19");
	mem(1152) := To_stdlogicvector(X"01");
	mem(1153) := To_stdlogicvector(X"13");
	mem(1154) := To_stdlogicvector(X"E0");
	mem(1155) := To_stdlogicvector(X"5F");
	mem(1156) := To_stdlogicvector(X"A0");
	mem(1157) := To_stdlogicvector(X"5D");
	mem(1158) := To_stdlogicvector(X"60");
	mem(1159) := To_stdlogicvector(X"5B");
	mem(1160) := To_stdlogicvector(X"20");
	mem(1161) := To_stdlogicvector(X"59");
	mem(1162) := To_stdlogicvector(X"0C");
	mem(1163) := To_stdlogicvector(X"64");
	mem(1164) := To_stdlogicvector(X"40");
	mem(1165) := To_stdlogicvector(X"66");
	mem(1166) := To_stdlogicvector(X"C4");
	mem(1167) := To_stdlogicvector(X"18");
	mem(1168) := To_stdlogicvector(X"62");
	mem(1169) := To_stdlogicvector(X"12");
	mem(1170) := To_stdlogicvector(X"BF");
	mem(1171) := To_stdlogicvector(X"14");
	mem(1172) := To_stdlogicvector(X"FB");
	mem(1173) := To_stdlogicvector(X"07");
	mem(1174) := To_stdlogicvector(X"22");
	mem(1175) := To_stdlogicvector(X"D9");
	mem(1176) := To_stdlogicvector(X"0C");
	mem(1177) := To_stdlogicvector(X"64");
	mem(1178) := To_stdlogicvector(X"40");
	mem(1179) := To_stdlogicvector(X"66");
	mem(1180) := To_stdlogicvector(X"C5");
	mem(1181) := To_stdlogicvector(X"1A");
	mem(1182) := To_stdlogicvector(X"62");
	mem(1183) := To_stdlogicvector(X"12");
	mem(1184) := To_stdlogicvector(X"BF");
	mem(1185) := To_stdlogicvector(X"14");
	mem(1186) := To_stdlogicvector(X"FB");
	mem(1187) := To_stdlogicvector(X"07");
	mem(1188) := To_stdlogicvector(X"62");
	mem(1189) := To_stdlogicvector(X"DB");
	mem(1190) := To_stdlogicvector(X"0C");
	mem(1191) := To_stdlogicvector(X"64");
	mem(1192) := To_stdlogicvector(X"40");
	mem(1193) := To_stdlogicvector(X"66");
	mem(1194) := To_stdlogicvector(X"C6");
	mem(1195) := To_stdlogicvector(X"1C");
	mem(1196) := To_stdlogicvector(X"62");
	mem(1197) := To_stdlogicvector(X"12");
	mem(1198) := To_stdlogicvector(X"BF");
	mem(1199) := To_stdlogicvector(X"14");
	mem(1200) := To_stdlogicvector(X"FB");
	mem(1201) := To_stdlogicvector(X"07");
	mem(1202) := To_stdlogicvector(X"A2");
	mem(1203) := To_stdlogicvector(X"DD");
	mem(1204) := To_stdlogicvector(X"0C");
	mem(1205) := To_stdlogicvector(X"64");
	mem(1206) := To_stdlogicvector(X"40");
	mem(1207) := To_stdlogicvector(X"66");
	mem(1208) := To_stdlogicvector(X"C7");
	mem(1209) := To_stdlogicvector(X"1E");
	mem(1210) := To_stdlogicvector(X"62");
	mem(1211) := To_stdlogicvector(X"12");
	mem(1212) := To_stdlogicvector(X"BF");
	mem(1213) := To_stdlogicvector(X"14");
	mem(1214) := To_stdlogicvector(X"FB");
	mem(1215) := To_stdlogicvector(X"07");
	mem(1216) := To_stdlogicvector(X"C7");
	mem(1217) := To_stdlogicvector(X"56");
	mem(1218) := To_stdlogicvector(X"FF");
	mem(1219) := To_stdlogicvector(X"9F");
	mem(1220) := To_stdlogicvector(X"FF");
	mem(1221) := To_stdlogicvector(X"0F");
	mem(1222) := To_stdlogicvector(X"00");
	mem(1223) := To_stdlogicvector(X"00");
	mem(1224) := To_stdlogicvector(X"00");
	mem(1225) := To_stdlogicvector(X"00");
	mem(1226) := To_stdlogicvector(X"00");
	mem(1227) := To_stdlogicvector(X"00");
	mem(1228) := To_stdlogicvector(X"00");
	mem(1229) := To_stdlogicvector(X"00");
	mem(1230) := To_stdlogicvector(X"00");
	mem(1231) := To_stdlogicvector(X"00");
	mem(1232) := To_stdlogicvector(X"00");
	mem(1233) := To_stdlogicvector(X"00");
	mem(1234) := To_stdlogicvector(X"00");
	mem(1235) := To_stdlogicvector(X"00");
	mem(1236) := To_stdlogicvector(X"00");
	mem(1237) := To_stdlogicvector(X"00");
	mem(1238) := To_stdlogicvector(X"00");
	mem(1239) := To_stdlogicvector(X"01");
	mem(1240) := To_stdlogicvector(X"00");
	mem(1241) := To_stdlogicvector(X"F0");
	mem(1242) := To_stdlogicvector(X"FF");
	mem(1243) := To_stdlogicvector(X"0F");
	mem(1244) := To_stdlogicvector(X"3F");
	mem(1245) := To_stdlogicvector(X"4A");
	mem(1246) := To_stdlogicvector(X"3F");
	mem(1247) := To_stdlogicvector(X"00");
	mem(1248) := To_stdlogicvector(X"F1");
	mem(1249) := To_stdlogicvector(X"FF");
	mem(1250) := To_stdlogicvector(X"FF");
	mem(1251) := To_stdlogicvector(X"00");
	mem(1252) := To_stdlogicvector(X"00");
	mem(1253) := To_stdlogicvector(X"00");
	mem(1254) := To_stdlogicvector(X"00");
	mem(1255) := To_stdlogicvector(X"00");
	mem(1256) := To_stdlogicvector(X"00");
	mem(1257) := To_stdlogicvector(X"00");
	mem(1258) := To_stdlogicvector(X"00");
	mem(1259) := To_stdlogicvector(X"00");
	mem(1260) := To_stdlogicvector(X"00");
	mem(1261) := To_stdlogicvector(X"00");
	mem(1262) := To_stdlogicvector(X"00");
	mem(1263) := To_stdlogicvector(X"00");
	mem(1264) := To_stdlogicvector(X"00");
	mem(1265) := To_stdlogicvector(X"00");
	mem(1266) := To_stdlogicvector(X"00");
	mem(1267) := To_stdlogicvector(X"00");
	mem(1268) := To_stdlogicvector(X"00");
	mem(1269) := To_stdlogicvector(X"00");
	mem(1270) := To_stdlogicvector(X"00");
	mem(1271) := To_stdlogicvector(X"00");
	mem(1272) := To_stdlogicvector(X"00");
	mem(1273) := To_stdlogicvector(X"00");
	mem(1274) := To_stdlogicvector(X"00");
	mem(1275) := To_stdlogicvector(X"00");
	mem(1276) := To_stdlogicvector(X"00");
	mem(1277) := To_stdlogicvector(X"00");
	mem(1278) := To_stdlogicvector(X"00");
	mem(1279) := To_stdlogicvector(X"00");
	mem(1280) := To_stdlogicvector(X"00");
	mem(1281) := To_stdlogicvector(X"00");
	mem(1282) := To_stdlogicvector(X"00");
	mem(1283) := To_stdlogicvector(X"00");
	mem(1284) := To_stdlogicvector(X"00");
	mem(1285) := To_stdlogicvector(X"00");
	mem(1286) := To_stdlogicvector(X"00");
	mem(1287) := To_stdlogicvector(X"00");
	mem(1288) := To_stdlogicvector(X"00");
	mem(1289) := To_stdlogicvector(X"00");
	mem(1290) := To_stdlogicvector(X"00");
	mem(1291) := To_stdlogicvector(X"00");
	mem(1292) := To_stdlogicvector(X"00");
	mem(1293) := To_stdlogicvector(X"00");
	mem(1294) := To_stdlogicvector(X"00");
	mem(1295) := To_stdlogicvector(X"00");
	mem(1296) := To_stdlogicvector(X"00");
	mem(1297) := To_stdlogicvector(X"00");
	mem(1298) := To_stdlogicvector(X"00");
	mem(1299) := To_stdlogicvector(X"00");
	mem(1300) := To_stdlogicvector(X"00");
	mem(1301) := To_stdlogicvector(X"00");
	mem(1302) := To_stdlogicvector(X"00");
	mem(1303) := To_stdlogicvector(X"00");
	mem(1304) := To_stdlogicvector(X"00");
	mem(1305) := To_stdlogicvector(X"00");
	mem(1306) := To_stdlogicvector(X"00");
	mem(1307) := To_stdlogicvector(X"00");
	mem(1308) := To_stdlogicvector(X"00");
	mem(1309) := To_stdlogicvector(X"00");
	mem(1310) := To_stdlogicvector(X"00");
	mem(1311) := To_stdlogicvector(X"00");
	mem(1312) := To_stdlogicvector(X"00");
	mem(1313) := To_stdlogicvector(X"00");
	mem(1314) := To_stdlogicvector(X"00");
	mem(1315) := To_stdlogicvector(X"00");
	mem(1316) := To_stdlogicvector(X"00");
	mem(1317) := To_stdlogicvector(X"00");
	mem(1318) := To_stdlogicvector(X"00");
	mem(1319) := To_stdlogicvector(X"00");
	mem(1320) := To_stdlogicvector(X"00");
	mem(1321) := To_stdlogicvector(X"00");
	mem(1322) := To_stdlogicvector(X"00");
	mem(1323) := To_stdlogicvector(X"00");
	mem(1324) := To_stdlogicvector(X"00");
	mem(1325) := To_stdlogicvector(X"00");
	mem(1326) := To_stdlogicvector(X"00");
	mem(1327) := To_stdlogicvector(X"00");
	mem(1328) := To_stdlogicvector(X"00");
	mem(1329) := To_stdlogicvector(X"00");
	mem(1330) := To_stdlogicvector(X"00");
	mem(1331) := To_stdlogicvector(X"00");
	mem(1332) := To_stdlogicvector(X"00");
	mem(1333) := To_stdlogicvector(X"00");
	mem(1334) := To_stdlogicvector(X"00");
	mem(1335) := To_stdlogicvector(X"00");
	mem(1336) := To_stdlogicvector(X"00");
	mem(1337) := To_stdlogicvector(X"00");
	mem(1338) := To_stdlogicvector(X"00");
	mem(1339) := To_stdlogicvector(X"00");
	mem(1340) := To_stdlogicvector(X"00");
	mem(1341) := To_stdlogicvector(X"00");
	mem(1342) := To_stdlogicvector(X"00");
	mem(1343) := To_stdlogicvector(X"00");
	mem(1344) := To_stdlogicvector(X"00");
	mem(1345) := To_stdlogicvector(X"00");
	mem(1346) := To_stdlogicvector(X"00");
	mem(1347) := To_stdlogicvector(X"00");
	mem(1348) := To_stdlogicvector(X"00");
	mem(1349) := To_stdlogicvector(X"00");
	mem(1350) := To_stdlogicvector(X"00");
	mem(1351) := To_stdlogicvector(X"00");
	mem(1352) := To_stdlogicvector(X"00");
	mem(1353) := To_stdlogicvector(X"00");
	mem(1354) := To_stdlogicvector(X"00");
	mem(1355) := To_stdlogicvector(X"00");
	mem(1356) := To_stdlogicvector(X"00");
	mem(1357) := To_stdlogicvector(X"00");
	mem(1358) := To_stdlogicvector(X"00");
	mem(1359) := To_stdlogicvector(X"00");
	mem(1360) := To_stdlogicvector(X"00");
	mem(1361) := To_stdlogicvector(X"00");
	mem(1362) := To_stdlogicvector(X"00");
	mem(1363) := To_stdlogicvector(X"00");
	mem(1364) := To_stdlogicvector(X"00");
	mem(1365) := To_stdlogicvector(X"00");
	mem(1366) := To_stdlogicvector(X"00");
	mem(1367) := To_stdlogicvector(X"00");
	mem(1368) := To_stdlogicvector(X"00");
	mem(1369) := To_stdlogicvector(X"00");
	mem(1370) := To_stdlogicvector(X"00");
	mem(1371) := To_stdlogicvector(X"00");
	mem(1372) := To_stdlogicvector(X"00");
	mem(1373) := To_stdlogicvector(X"00");
	mem(1374) := To_stdlogicvector(X"00");
	mem(1375) := To_stdlogicvector(X"00");
	mem(1376) := To_stdlogicvector(X"00");
	mem(1377) := To_stdlogicvector(X"00");
	mem(1378) := To_stdlogicvector(X"00");
	mem(1379) := To_stdlogicvector(X"00");
	mem(1380) := To_stdlogicvector(X"00");
	mem(1381) := To_stdlogicvector(X"00");
	mem(1382) := To_stdlogicvector(X"00");
	mem(1383) := To_stdlogicvector(X"00");
	mem(1384) := To_stdlogicvector(X"00");
	mem(1385) := To_stdlogicvector(X"00");
	mem(1386) := To_stdlogicvector(X"00");
	mem(1387) := To_stdlogicvector(X"00");
	mem(1388) := To_stdlogicvector(X"00");
	mem(1389) := To_stdlogicvector(X"00");
	mem(1390) := To_stdlogicvector(X"00");
	mem(1391) := To_stdlogicvector(X"00");
	mem(1392) := To_stdlogicvector(X"00");
	mem(1393) := To_stdlogicvector(X"00");
	mem(1394) := To_stdlogicvector(X"00");
	mem(1395) := To_stdlogicvector(X"00");
	mem(1396) := To_stdlogicvector(X"00");
	mem(1397) := To_stdlogicvector(X"00");
	mem(1398) := To_stdlogicvector(X"00");
	mem(1399) := To_stdlogicvector(X"00");
	mem(1400) := To_stdlogicvector(X"00");
	mem(1401) := To_stdlogicvector(X"00");
	mem(1402) := To_stdlogicvector(X"00");
	mem(1403) := To_stdlogicvector(X"00");
	mem(1404) := To_stdlogicvector(X"00");
	mem(1405) := To_stdlogicvector(X"00");
	mem(1406) := To_stdlogicvector(X"00");
	mem(1407) := To_stdlogicvector(X"00");
	mem(1408) := To_stdlogicvector(X"00");
	mem(1409) := To_stdlogicvector(X"00");
	mem(1410) := To_stdlogicvector(X"00");
	mem(1411) := To_stdlogicvector(X"00");
	mem(1412) := To_stdlogicvector(X"00");
	mem(1413) := To_stdlogicvector(X"00");
	mem(1414) := To_stdlogicvector(X"00");
	mem(1415) := To_stdlogicvector(X"00");
	mem(1416) := To_stdlogicvector(X"00");
	mem(1417) := To_stdlogicvector(X"00");
	mem(1418) := To_stdlogicvector(X"00");
	mem(1419) := To_stdlogicvector(X"00");
	mem(1420) := To_stdlogicvector(X"00");
	mem(1421) := To_stdlogicvector(X"00");
	mem(1422) := To_stdlogicvector(X"00");
	mem(1423) := To_stdlogicvector(X"00");
	mem(1424) := To_stdlogicvector(X"00");
	mem(1425) := To_stdlogicvector(X"00");
	mem(1426) := To_stdlogicvector(X"00");
	mem(1427) := To_stdlogicvector(X"00");
	mem(1428) := To_stdlogicvector(X"00");
	mem(1429) := To_stdlogicvector(X"00");
	mem(1430) := To_stdlogicvector(X"00");
	mem(1431) := To_stdlogicvector(X"00");
	mem(1432) := To_stdlogicvector(X"00");
	mem(1433) := To_stdlogicvector(X"00");
	mem(1434) := To_stdlogicvector(X"00");
	mem(1435) := To_stdlogicvector(X"00");
	mem(1436) := To_stdlogicvector(X"00");
	mem(1437) := To_stdlogicvector(X"00");
	mem(1438) := To_stdlogicvector(X"00");
	mem(1439) := To_stdlogicvector(X"00");
	mem(1440) := To_stdlogicvector(X"00");
	mem(1441) := To_stdlogicvector(X"00");
	mem(1442) := To_stdlogicvector(X"00");
	mem(1443) := To_stdlogicvector(X"00");
	mem(1444) := To_stdlogicvector(X"00");
	mem(1445) := To_stdlogicvector(X"00");
	mem(1446) := To_stdlogicvector(X"00");
	mem(1447) := To_stdlogicvector(X"00");
	mem(1448) := To_stdlogicvector(X"00");
	mem(1449) := To_stdlogicvector(X"00");
	mem(1450) := To_stdlogicvector(X"00");
	mem(1451) := To_stdlogicvector(X"00");
	mem(1452) := To_stdlogicvector(X"00");
	mem(1453) := To_stdlogicvector(X"00");
	mem(1454) := To_stdlogicvector(X"00");
	mem(1455) := To_stdlogicvector(X"00");
	mem(1456) := To_stdlogicvector(X"00");
	mem(1457) := To_stdlogicvector(X"00");
	mem(1458) := To_stdlogicvector(X"00");
	mem(1459) := To_stdlogicvector(X"00");
	mem(1460) := To_stdlogicvector(X"00");
	mem(1461) := To_stdlogicvector(X"00");
	mem(1462) := To_stdlogicvector(X"00");
	mem(1463) := To_stdlogicvector(X"00");
	mem(1464) := To_stdlogicvector(X"00");
	mem(1465) := To_stdlogicvector(X"00");
	mem(1466) := To_stdlogicvector(X"00");
	mem(1467) := To_stdlogicvector(X"00");
	mem(1468) := To_stdlogicvector(X"00");
	mem(1469) := To_stdlogicvector(X"00");
	mem(1470) := To_stdlogicvector(X"00");
	mem(1471) := To_stdlogicvector(X"00");
	mem(1472) := To_stdlogicvector(X"00");
	mem(1473) := To_stdlogicvector(X"00");
	mem(1474) := To_stdlogicvector(X"00");
	mem(1475) := To_stdlogicvector(X"00");
	mem(1476) := To_stdlogicvector(X"00");
	mem(1477) := To_stdlogicvector(X"00");
	mem(1478) := To_stdlogicvector(X"00");
	mem(1479) := To_stdlogicvector(X"00");
	mem(1480) := To_stdlogicvector(X"00");
	mem(1481) := To_stdlogicvector(X"00");
	mem(1482) := To_stdlogicvector(X"00");
	mem(1483) := To_stdlogicvector(X"00");
	mem(1484) := To_stdlogicvector(X"00");
	mem(1485) := To_stdlogicvector(X"00");
	mem(1486) := To_stdlogicvector(X"00");
	mem(1487) := To_stdlogicvector(X"00");
	mem(1488) := To_stdlogicvector(X"00");
	mem(1489) := To_stdlogicvector(X"00");
	mem(1490) := To_stdlogicvector(X"00");
	mem(1491) := To_stdlogicvector(X"00");
	mem(1492) := To_stdlogicvector(X"00");
	mem(1493) := To_stdlogicvector(X"00");
	mem(1494) := To_stdlogicvector(X"00");
	mem(1495) := To_stdlogicvector(X"00");
	mem(1496) := To_stdlogicvector(X"00");
	mem(1497) := To_stdlogicvector(X"00");
	mem(1498) := To_stdlogicvector(X"00");
	mem(1499) := To_stdlogicvector(X"00");
	mem(1500) := To_stdlogicvector(X"00");
	mem(1501) := To_stdlogicvector(X"00");
	mem(1502) := To_stdlogicvector(X"00");
	mem(1503) := To_stdlogicvector(X"00");
	mem(1504) := To_stdlogicvector(X"00");
	mem(1505) := To_stdlogicvector(X"00");
	mem(1506) := To_stdlogicvector(X"00");
	mem(1507) := To_stdlogicvector(X"00");
	mem(1508) := To_stdlogicvector(X"00");
	mem(1509) := To_stdlogicvector(X"00");
	mem(1510) := To_stdlogicvector(X"00");
	mem(1511) := To_stdlogicvector(X"00");
	mem(1512) := To_stdlogicvector(X"00");
	mem(1513) := To_stdlogicvector(X"00");
	mem(1514) := To_stdlogicvector(X"00");
	mem(1515) := To_stdlogicvector(X"00");
	mem(1516) := To_stdlogicvector(X"00");
	mem(1517) := To_stdlogicvector(X"00");
	mem(1518) := To_stdlogicvector(X"00");
	mem(1519) := To_stdlogicvector(X"00");
	mem(1520) := To_stdlogicvector(X"00");
	mem(1521) := To_stdlogicvector(X"00");
	mem(1522) := To_stdlogicvector(X"00");
	mem(1523) := To_stdlogicvector(X"00");
	mem(1524) := To_stdlogicvector(X"00");
	mem(1525) := To_stdlogicvector(X"00");
	mem(1526) := To_stdlogicvector(X"00");
	mem(1527) := To_stdlogicvector(X"00");
	mem(1528) := To_stdlogicvector(X"00");
	mem(1529) := To_stdlogicvector(X"00");
	mem(1530) := To_stdlogicvector(X"00");
	mem(1531) := To_stdlogicvector(X"00");
	mem(1532) := To_stdlogicvector(X"00");
	mem(1533) := To_stdlogicvector(X"00");
	mem(1534) := To_stdlogicvector(X"00");
	mem(1535) := To_stdlogicvector(X"00");
	mem(1536) := To_stdlogicvector(X"00");
	mem(1537) := To_stdlogicvector(X"00");
	mem(1538) := To_stdlogicvector(X"00");
	mem(1539) := To_stdlogicvector(X"00");
	mem(1540) := To_stdlogicvector(X"00");
	mem(1541) := To_stdlogicvector(X"00");
	mem(1542) := To_stdlogicvector(X"00");
	mem(1543) := To_stdlogicvector(X"00");
	mem(1544) := To_stdlogicvector(X"00");
	mem(1545) := To_stdlogicvector(X"00");
	mem(1546) := To_stdlogicvector(X"00");
	mem(1547) := To_stdlogicvector(X"00");
	mem(1548) := To_stdlogicvector(X"00");
	mem(1549) := To_stdlogicvector(X"00");
	mem(1550) := To_stdlogicvector(X"00");
	mem(1551) := To_stdlogicvector(X"00");
	mem(1552) := To_stdlogicvector(X"00");
	mem(1553) := To_stdlogicvector(X"00");
	mem(1554) := To_stdlogicvector(X"00");
	mem(1555) := To_stdlogicvector(X"00");
	mem(1556) := To_stdlogicvector(X"00");
	mem(1557) := To_stdlogicvector(X"00");
	mem(1558) := To_stdlogicvector(X"00");
	mem(1559) := To_stdlogicvector(X"00");
	mem(1560) := To_stdlogicvector(X"00");
	mem(1561) := To_stdlogicvector(X"00");
	mem(1562) := To_stdlogicvector(X"00");
	mem(1563) := To_stdlogicvector(X"00");
	mem(1564) := To_stdlogicvector(X"00");
	mem(1565) := To_stdlogicvector(X"00");
	mem(1566) := To_stdlogicvector(X"00");
	mem(1567) := To_stdlogicvector(X"00");
	mem(1568) := To_stdlogicvector(X"00");
	mem(1569) := To_stdlogicvector(X"00");
	mem(1570) := To_stdlogicvector(X"00");
	mem(1571) := To_stdlogicvector(X"00");
	mem(1572) := To_stdlogicvector(X"00");
	mem(1573) := To_stdlogicvector(X"00");
	mem(1574) := To_stdlogicvector(X"00");
	mem(1575) := To_stdlogicvector(X"00");
	mem(1576) := To_stdlogicvector(X"00");
	mem(1577) := To_stdlogicvector(X"00");
	mem(1578) := To_stdlogicvector(X"00");
	mem(1579) := To_stdlogicvector(X"00");
	mem(1580) := To_stdlogicvector(X"00");
	mem(1581) := To_stdlogicvector(X"00");
	mem(1582) := To_stdlogicvector(X"00");
	mem(1583) := To_stdlogicvector(X"00");
	mem(1584) := To_stdlogicvector(X"00");
	mem(1585) := To_stdlogicvector(X"00");
	mem(1586) := To_stdlogicvector(X"00");
	mem(1587) := To_stdlogicvector(X"00");
	mem(1588) := To_stdlogicvector(X"00");
	mem(1589) := To_stdlogicvector(X"00");
	mem(1590) := To_stdlogicvector(X"00");
	mem(1591) := To_stdlogicvector(X"00");
	mem(1592) := To_stdlogicvector(X"00");
	mem(1593) := To_stdlogicvector(X"00");
	mem(1594) := To_stdlogicvector(X"00");
	mem(1595) := To_stdlogicvector(X"00");
	mem(1596) := To_stdlogicvector(X"00");
	mem(1597) := To_stdlogicvector(X"00");
	mem(1598) := To_stdlogicvector(X"00");
	mem(1599) := To_stdlogicvector(X"00");
	mem(1600) := To_stdlogicvector(X"00");
	mem(1601) := To_stdlogicvector(X"00");
	mem(1602) := To_stdlogicvector(X"00");
	mem(1603) := To_stdlogicvector(X"00");
	mem(1604) := To_stdlogicvector(X"00");
	mem(1605) := To_stdlogicvector(X"00");
	mem(1606) := To_stdlogicvector(X"00");
	mem(1607) := To_stdlogicvector(X"00");
	mem(1608) := To_stdlogicvector(X"00");
	mem(1609) := To_stdlogicvector(X"00");
	mem(1610) := To_stdlogicvector(X"00");
	mem(1611) := To_stdlogicvector(X"00");
	mem(1612) := To_stdlogicvector(X"00");
	mem(1613) := To_stdlogicvector(X"00");
	mem(1614) := To_stdlogicvector(X"00");
	mem(1615) := To_stdlogicvector(X"00");
	mem(1616) := To_stdlogicvector(X"00");
	mem(1617) := To_stdlogicvector(X"00");
	mem(1618) := To_stdlogicvector(X"00");
	mem(1619) := To_stdlogicvector(X"00");
	mem(1620) := To_stdlogicvector(X"00");
	mem(1621) := To_stdlogicvector(X"00");
	mem(1622) := To_stdlogicvector(X"00");
	mem(1623) := To_stdlogicvector(X"00");
	mem(1624) := To_stdlogicvector(X"00");
	mem(1625) := To_stdlogicvector(X"00");
	mem(1626) := To_stdlogicvector(X"00");
	mem(1627) := To_stdlogicvector(X"00");
	mem(1628) := To_stdlogicvector(X"00");
	mem(1629) := To_stdlogicvector(X"00");
	mem(1630) := To_stdlogicvector(X"00");
	mem(1631) := To_stdlogicvector(X"00");
	mem(1632) := To_stdlogicvector(X"00");
	mem(1633) := To_stdlogicvector(X"00");
	mem(1634) := To_stdlogicvector(X"00");
	mem(1635) := To_stdlogicvector(X"00");
	mem(1636) := To_stdlogicvector(X"00");
	mem(1637) := To_stdlogicvector(X"00");
	mem(1638) := To_stdlogicvector(X"00");
	mem(1639) := To_stdlogicvector(X"00");
	mem(1640) := To_stdlogicvector(X"00");
	mem(1641) := To_stdlogicvector(X"00");
	mem(1642) := To_stdlogicvector(X"00");
	mem(1643) := To_stdlogicvector(X"00");
	mem(1644) := To_stdlogicvector(X"00");
	mem(1645) := To_stdlogicvector(X"00");
	mem(1646) := To_stdlogicvector(X"00");
	mem(1647) := To_stdlogicvector(X"00");
	mem(1648) := To_stdlogicvector(X"00");
	mem(1649) := To_stdlogicvector(X"00");
	mem(1650) := To_stdlogicvector(X"00");
	mem(1651) := To_stdlogicvector(X"00");
	mem(1652) := To_stdlogicvector(X"00");
	mem(1653) := To_stdlogicvector(X"00");
	mem(1654) := To_stdlogicvector(X"00");
	mem(1655) := To_stdlogicvector(X"00");
	mem(1656) := To_stdlogicvector(X"00");
	mem(1657) := To_stdlogicvector(X"00");
	mem(1658) := To_stdlogicvector(X"00");
	mem(1659) := To_stdlogicvector(X"00");
	mem(1660) := To_stdlogicvector(X"00");
	mem(1661) := To_stdlogicvector(X"00");
	mem(1662) := To_stdlogicvector(X"00");
	mem(1663) := To_stdlogicvector(X"00");
	mem(1664) := To_stdlogicvector(X"00");
	mem(1665) := To_stdlogicvector(X"00");
	mem(1666) := To_stdlogicvector(X"00");
	mem(1667) := To_stdlogicvector(X"00");
	mem(1668) := To_stdlogicvector(X"00");
	mem(1669) := To_stdlogicvector(X"00");
	mem(1670) := To_stdlogicvector(X"00");
	mem(1671) := To_stdlogicvector(X"00");
	mem(1672) := To_stdlogicvector(X"00");
	mem(1673) := To_stdlogicvector(X"00");
	mem(1674) := To_stdlogicvector(X"00");
	mem(1675) := To_stdlogicvector(X"00");
	mem(1676) := To_stdlogicvector(X"00");
	mem(1677) := To_stdlogicvector(X"00");
	mem(1678) := To_stdlogicvector(X"00");
	mem(1679) := To_stdlogicvector(X"00");
	mem(1680) := To_stdlogicvector(X"00");
	mem(1681) := To_stdlogicvector(X"00");
	mem(1682) := To_stdlogicvector(X"00");
	mem(1683) := To_stdlogicvector(X"00");
	mem(1684) := To_stdlogicvector(X"00");
	mem(1685) := To_stdlogicvector(X"00");
	mem(1686) := To_stdlogicvector(X"00");
	mem(1687) := To_stdlogicvector(X"00");
	mem(1688) := To_stdlogicvector(X"00");
	mem(1689) := To_stdlogicvector(X"00");
	mem(1690) := To_stdlogicvector(X"00");
	mem(1691) := To_stdlogicvector(X"00");
	mem(1692) := To_stdlogicvector(X"00");
	mem(1693) := To_stdlogicvector(X"00");
	mem(1694) := To_stdlogicvector(X"00");
	mem(1695) := To_stdlogicvector(X"00");
	mem(1696) := To_stdlogicvector(X"00");
	mem(1697) := To_stdlogicvector(X"00");
	mem(1698) := To_stdlogicvector(X"00");
	mem(1699) := To_stdlogicvector(X"00");
	mem(1700) := To_stdlogicvector(X"00");
	mem(1701) := To_stdlogicvector(X"00");
	mem(1702) := To_stdlogicvector(X"00");
	mem(1703) := To_stdlogicvector(X"00");
	mem(1704) := To_stdlogicvector(X"00");
	mem(1705) := To_stdlogicvector(X"00");
	mem(1706) := To_stdlogicvector(X"00");
	mem(1707) := To_stdlogicvector(X"00");
	mem(1708) := To_stdlogicvector(X"00");
	mem(1709) := To_stdlogicvector(X"00");
	mem(1710) := To_stdlogicvector(X"00");
	mem(1711) := To_stdlogicvector(X"00");
	mem(1712) := To_stdlogicvector(X"00");
	mem(1713) := To_stdlogicvector(X"00");
	mem(1714) := To_stdlogicvector(X"00");
	mem(1715) := To_stdlogicvector(X"00");
	mem(1716) := To_stdlogicvector(X"00");
	mem(1717) := To_stdlogicvector(X"00");
	mem(1718) := To_stdlogicvector(X"00");
	mem(1719) := To_stdlogicvector(X"00");
	mem(1720) := To_stdlogicvector(X"00");
	mem(1721) := To_stdlogicvector(X"00");
	mem(1722) := To_stdlogicvector(X"00");
	mem(1723) := To_stdlogicvector(X"00");
	mem(1724) := To_stdlogicvector(X"00");
	mem(1725) := To_stdlogicvector(X"00");
	mem(1726) := To_stdlogicvector(X"00");
	mem(1727) := To_stdlogicvector(X"00");
	mem(1728) := To_stdlogicvector(X"00");
	mem(1729) := To_stdlogicvector(X"00");
	mem(1730) := To_stdlogicvector(X"00");
	mem(1731) := To_stdlogicvector(X"00");
	mem(1732) := To_stdlogicvector(X"00");
	mem(1733) := To_stdlogicvector(X"00");
	mem(1734) := To_stdlogicvector(X"00");
	mem(1735) := To_stdlogicvector(X"00");
	mem(1736) := To_stdlogicvector(X"00");
	mem(1737) := To_stdlogicvector(X"00");
	mem(1738) := To_stdlogicvector(X"00");
	mem(1739) := To_stdlogicvector(X"00");
	mem(1740) := To_stdlogicvector(X"00");
	mem(1741) := To_stdlogicvector(X"00");
	mem(1742) := To_stdlogicvector(X"00");
	mem(1743) := To_stdlogicvector(X"00");
	mem(1744) := To_stdlogicvector(X"00");
	mem(1745) := To_stdlogicvector(X"00");
	mem(1746) := To_stdlogicvector(X"00");
	mem(1747) := To_stdlogicvector(X"00");
	mem(1748) := To_stdlogicvector(X"00");
	mem(1749) := To_stdlogicvector(X"00");
	mem(1750) := To_stdlogicvector(X"00");
	mem(1751) := To_stdlogicvector(X"00");
	mem(1752) := To_stdlogicvector(X"00");
	mem(1753) := To_stdlogicvector(X"00");
	mem(1754) := To_stdlogicvector(X"00");
	mem(1755) := To_stdlogicvector(X"00");
	mem(1756) := To_stdlogicvector(X"00");
	mem(1757) := To_stdlogicvector(X"00");
	mem(1758) := To_stdlogicvector(X"00");
	mem(1759) := To_stdlogicvector(X"00");
	mem(1760) := To_stdlogicvector(X"00");
	mem(1761) := To_stdlogicvector(X"00");
	mem(1762) := To_stdlogicvector(X"00");
	mem(1763) := To_stdlogicvector(X"00");
	mem(1764) := To_stdlogicvector(X"00");
	mem(1765) := To_stdlogicvector(X"00");
	mem(1766) := To_stdlogicvector(X"00");
	mem(1767) := To_stdlogicvector(X"00");
	mem(1768) := To_stdlogicvector(X"00");
	mem(1769) := To_stdlogicvector(X"00");
	mem(1770) := To_stdlogicvector(X"00");
	mem(1771) := To_stdlogicvector(X"00");
	mem(1772) := To_stdlogicvector(X"00");
	mem(1773) := To_stdlogicvector(X"00");
	mem(1774) := To_stdlogicvector(X"00");
	mem(1775) := To_stdlogicvector(X"00");
	mem(1776) := To_stdlogicvector(X"00");
	mem(1777) := To_stdlogicvector(X"00");
	mem(1778) := To_stdlogicvector(X"00");
	mem(1779) := To_stdlogicvector(X"00");
	mem(1780) := To_stdlogicvector(X"00");
	mem(1781) := To_stdlogicvector(X"00");
	mem(1782) := To_stdlogicvector(X"00");
	mem(1783) := To_stdlogicvector(X"00");
	mem(1784) := To_stdlogicvector(X"00");
	mem(1785) := To_stdlogicvector(X"00");
	mem(1786) := To_stdlogicvector(X"00");
	mem(1787) := To_stdlogicvector(X"00");
	mem(1788) := To_stdlogicvector(X"00");
	mem(1789) := To_stdlogicvector(X"00");
	mem(1790) := To_stdlogicvector(X"00");
	mem(1791) := To_stdlogicvector(X"00");
	mem(1792) := To_stdlogicvector(X"00");
	mem(1793) := To_stdlogicvector(X"00");
	mem(1794) := To_stdlogicvector(X"00");
	mem(1795) := To_stdlogicvector(X"00");
	mem(1796) := To_stdlogicvector(X"00");
	mem(1797) := To_stdlogicvector(X"00");
	mem(1798) := To_stdlogicvector(X"00");
	mem(1799) := To_stdlogicvector(X"00");
	mem(1800) := To_stdlogicvector(X"00");
	mem(1801) := To_stdlogicvector(X"00");
	mem(1802) := To_stdlogicvector(X"00");
	mem(1803) := To_stdlogicvector(X"00");
	mem(1804) := To_stdlogicvector(X"00");
	mem(1805) := To_stdlogicvector(X"00");
	mem(1806) := To_stdlogicvector(X"00");
	mem(1807) := To_stdlogicvector(X"00");
	mem(1808) := To_stdlogicvector(X"00");
	mem(1809) := To_stdlogicvector(X"00");
	mem(1810) := To_stdlogicvector(X"00");
	mem(1811) := To_stdlogicvector(X"00");
	mem(1812) := To_stdlogicvector(X"00");
	mem(1813) := To_stdlogicvector(X"00");
	mem(1814) := To_stdlogicvector(X"00");
	mem(1815) := To_stdlogicvector(X"00");
	mem(1816) := To_stdlogicvector(X"00");
	mem(1817) := To_stdlogicvector(X"00");
	mem(1818) := To_stdlogicvector(X"00");
	mem(1819) := To_stdlogicvector(X"00");
	mem(1820) := To_stdlogicvector(X"00");
	mem(1821) := To_stdlogicvector(X"00");
	mem(1822) := To_stdlogicvector(X"00");
	mem(1823) := To_stdlogicvector(X"00");
	mem(1824) := To_stdlogicvector(X"00");
	mem(1825) := To_stdlogicvector(X"00");
	mem(1826) := To_stdlogicvector(X"00");
	mem(1827) := To_stdlogicvector(X"00");
	mem(1828) := To_stdlogicvector(X"00");
	mem(1829) := To_stdlogicvector(X"00");
	mem(1830) := To_stdlogicvector(X"00");
	mem(1831) := To_stdlogicvector(X"00");
	mem(1832) := To_stdlogicvector(X"00");
	mem(1833) := To_stdlogicvector(X"00");
	mem(1834) := To_stdlogicvector(X"00");
	mem(1835) := To_stdlogicvector(X"00");
	mem(1836) := To_stdlogicvector(X"00");
	mem(1837) := To_stdlogicvector(X"00");
	mem(1838) := To_stdlogicvector(X"00");
	mem(1839) := To_stdlogicvector(X"00");
	mem(1840) := To_stdlogicvector(X"00");
	mem(1841) := To_stdlogicvector(X"00");
	mem(1842) := To_stdlogicvector(X"00");
	mem(1843) := To_stdlogicvector(X"00");
	mem(1844) := To_stdlogicvector(X"00");
	mem(1845) := To_stdlogicvector(X"00");
	mem(1846) := To_stdlogicvector(X"00");
	mem(1847) := To_stdlogicvector(X"00");
	mem(1848) := To_stdlogicvector(X"00");
	mem(1849) := To_stdlogicvector(X"00");
	mem(1850) := To_stdlogicvector(X"00");
	mem(1851) := To_stdlogicvector(X"00");
	mem(1852) := To_stdlogicvector(X"00");
	mem(1853) := To_stdlogicvector(X"00");
	mem(1854) := To_stdlogicvector(X"00");
	mem(1855) := To_stdlogicvector(X"00");
	mem(1856) := To_stdlogicvector(X"00");
	mem(1857) := To_stdlogicvector(X"00");
	mem(1858) := To_stdlogicvector(X"00");
	mem(1859) := To_stdlogicvector(X"00");
	mem(1860) := To_stdlogicvector(X"00");
	mem(1861) := To_stdlogicvector(X"00");
	mem(1862) := To_stdlogicvector(X"00");
	mem(1863) := To_stdlogicvector(X"00");
	mem(1864) := To_stdlogicvector(X"00");
	mem(1865) := To_stdlogicvector(X"00");
	mem(1866) := To_stdlogicvector(X"00");
	mem(1867) := To_stdlogicvector(X"00");
	mem(1868) := To_stdlogicvector(X"00");
	mem(1869) := To_stdlogicvector(X"00");
	mem(1870) := To_stdlogicvector(X"00");
	mem(1871) := To_stdlogicvector(X"00");
	mem(1872) := To_stdlogicvector(X"00");
	mem(1873) := To_stdlogicvector(X"00");
	mem(1874) := To_stdlogicvector(X"00");
	mem(1875) := To_stdlogicvector(X"00");
	mem(1876) := To_stdlogicvector(X"00");
	mem(1877) := To_stdlogicvector(X"00");
	mem(1878) := To_stdlogicvector(X"00");
	mem(1879) := To_stdlogicvector(X"00");
	mem(1880) := To_stdlogicvector(X"00");
	mem(1881) := To_stdlogicvector(X"00");
	mem(1882) := To_stdlogicvector(X"00");
	mem(1883) := To_stdlogicvector(X"00");
	mem(1884) := To_stdlogicvector(X"00");
	mem(1885) := To_stdlogicvector(X"00");
	mem(1886) := To_stdlogicvector(X"00");
	mem(1887) := To_stdlogicvector(X"00");
	mem(1888) := To_stdlogicvector(X"00");
	mem(1889) := To_stdlogicvector(X"00");
	mem(1890) := To_stdlogicvector(X"00");
	mem(1891) := To_stdlogicvector(X"00");
	mem(1892) := To_stdlogicvector(X"00");
	mem(1893) := To_stdlogicvector(X"00");
	mem(1894) := To_stdlogicvector(X"00");
	mem(1895) := To_stdlogicvector(X"00");
	mem(1896) := To_stdlogicvector(X"00");
	mem(1897) := To_stdlogicvector(X"00");
	mem(1898) := To_stdlogicvector(X"00");
	mem(1899) := To_stdlogicvector(X"00");
	mem(1900) := To_stdlogicvector(X"00");
	mem(1901) := To_stdlogicvector(X"00");
	mem(1902) := To_stdlogicvector(X"00");
	mem(1903) := To_stdlogicvector(X"00");
	mem(1904) := To_stdlogicvector(X"00");
	mem(1905) := To_stdlogicvector(X"00");
	mem(1906) := To_stdlogicvector(X"00");
	mem(1907) := To_stdlogicvector(X"00");
	mem(1908) := To_stdlogicvector(X"00");
	mem(1909) := To_stdlogicvector(X"00");
	mem(1910) := To_stdlogicvector(X"00");
	mem(1911) := To_stdlogicvector(X"00");
	mem(1912) := To_stdlogicvector(X"00");
	mem(1913) := To_stdlogicvector(X"00");
	mem(1914) := To_stdlogicvector(X"00");
	mem(1915) := To_stdlogicvector(X"00");
	mem(1916) := To_stdlogicvector(X"00");
	mem(1917) := To_stdlogicvector(X"00");
	mem(1918) := To_stdlogicvector(X"00");
	mem(1919) := To_stdlogicvector(X"00");
	mem(1920) := To_stdlogicvector(X"00");
	mem(1921) := To_stdlogicvector(X"00");
	mem(1922) := To_stdlogicvector(X"00");
	mem(1923) := To_stdlogicvector(X"00");
	mem(1924) := To_stdlogicvector(X"00");
	mem(1925) := To_stdlogicvector(X"00");
	mem(1926) := To_stdlogicvector(X"00");
	mem(1927) := To_stdlogicvector(X"00");
	mem(1928) := To_stdlogicvector(X"00");
	mem(1929) := To_stdlogicvector(X"00");
	mem(1930) := To_stdlogicvector(X"00");
	mem(1931) := To_stdlogicvector(X"00");
	mem(1932) := To_stdlogicvector(X"00");
	mem(1933) := To_stdlogicvector(X"00");
	mem(1934) := To_stdlogicvector(X"00");
	mem(1935) := To_stdlogicvector(X"00");
	mem(1936) := To_stdlogicvector(X"00");
	mem(1937) := To_stdlogicvector(X"00");
	mem(1938) := To_stdlogicvector(X"00");
	mem(1939) := To_stdlogicvector(X"00");
	mem(1940) := To_stdlogicvector(X"00");
	mem(1941) := To_stdlogicvector(X"00");
	mem(1942) := To_stdlogicvector(X"00");
	mem(1943) := To_stdlogicvector(X"00");
	mem(1944) := To_stdlogicvector(X"00");
	mem(1945) := To_stdlogicvector(X"00");
	mem(1946) := To_stdlogicvector(X"00");
	mem(1947) := To_stdlogicvector(X"00");
	mem(1948) := To_stdlogicvector(X"00");
	mem(1949) := To_stdlogicvector(X"00");
	mem(1950) := To_stdlogicvector(X"00");
	mem(1951) := To_stdlogicvector(X"00");
	mem(1952) := To_stdlogicvector(X"00");
	mem(1953) := To_stdlogicvector(X"00");
	mem(1954) := To_stdlogicvector(X"00");
	mem(1955) := To_stdlogicvector(X"00");
	mem(1956) := To_stdlogicvector(X"00");
	mem(1957) := To_stdlogicvector(X"00");
	mem(1958) := To_stdlogicvector(X"00");
	mem(1959) := To_stdlogicvector(X"00");
	mem(1960) := To_stdlogicvector(X"00");
	mem(1961) := To_stdlogicvector(X"00");
	mem(1962) := To_stdlogicvector(X"00");
	mem(1963) := To_stdlogicvector(X"00");
	mem(1964) := To_stdlogicvector(X"00");
	mem(1965) := To_stdlogicvector(X"00");
	mem(1966) := To_stdlogicvector(X"00");
	mem(1967) := To_stdlogicvector(X"00");
	mem(1968) := To_stdlogicvector(X"00");
	mem(1969) := To_stdlogicvector(X"00");
	mem(1970) := To_stdlogicvector(X"00");
	mem(1971) := To_stdlogicvector(X"00");
	mem(1972) := To_stdlogicvector(X"00");
	mem(1973) := To_stdlogicvector(X"00");
	mem(1974) := To_stdlogicvector(X"00");
	mem(1975) := To_stdlogicvector(X"00");
	mem(1976) := To_stdlogicvector(X"00");
	mem(1977) := To_stdlogicvector(X"00");
	mem(1978) := To_stdlogicvector(X"00");
	mem(1979) := To_stdlogicvector(X"00");
	mem(1980) := To_stdlogicvector(X"00");
	mem(1981) := To_stdlogicvector(X"00");
	mem(1982) := To_stdlogicvector(X"00");
	mem(1983) := To_stdlogicvector(X"00");
	mem(1984) := To_stdlogicvector(X"00");
	mem(1985) := To_stdlogicvector(X"00");
	mem(1986) := To_stdlogicvector(X"00");
	mem(1987) := To_stdlogicvector(X"00");
	mem(1988) := To_stdlogicvector(X"00");
	mem(1989) := To_stdlogicvector(X"00");
	mem(1990) := To_stdlogicvector(X"00");
	mem(1991) := To_stdlogicvector(X"00");
	mem(1992) := To_stdlogicvector(X"00");
	mem(1993) := To_stdlogicvector(X"00");
	mem(1994) := To_stdlogicvector(X"00");
	mem(1995) := To_stdlogicvector(X"00");
	mem(1996) := To_stdlogicvector(X"00");
	mem(1997) := To_stdlogicvector(X"00");
	mem(1998) := To_stdlogicvector(X"00");
	mem(1999) := To_stdlogicvector(X"00");
	mem(2000) := To_stdlogicvector(X"00");
	mem(2001) := To_stdlogicvector(X"00");
	mem(2002) := To_stdlogicvector(X"00");
	mem(2003) := To_stdlogicvector(X"00");
	mem(2004) := To_stdlogicvector(X"00");
	mem(2005) := To_stdlogicvector(X"00");
	mem(2006) := To_stdlogicvector(X"00");
	mem(2007) := To_stdlogicvector(X"00");
	mem(2008) := To_stdlogicvector(X"00");
	mem(2009) := To_stdlogicvector(X"00");
	mem(2010) := To_stdlogicvector(X"00");
	mem(2011) := To_stdlogicvector(X"00");
	mem(2012) := To_stdlogicvector(X"00");
	mem(2013) := To_stdlogicvector(X"00");
	mem(2014) := To_stdlogicvector(X"00");
	mem(2015) := To_stdlogicvector(X"00");
	mem(2016) := To_stdlogicvector(X"00");
	mem(2017) := To_stdlogicvector(X"00");
	mem(2018) := To_stdlogicvector(X"00");
	mem(2019) := To_stdlogicvector(X"00");
	mem(2020) := To_stdlogicvector(X"00");
	mem(2021) := To_stdlogicvector(X"00");
	mem(2022) := To_stdlogicvector(X"00");
	mem(2023) := To_stdlogicvector(X"00");
	mem(2024) := To_stdlogicvector(X"00");
	mem(2025) := To_stdlogicvector(X"00");
	mem(2026) := To_stdlogicvector(X"00");
	mem(2027) := To_stdlogicvector(X"00");
	mem(2028) := To_stdlogicvector(X"00");
	mem(2029) := To_stdlogicvector(X"00");
	mem(2030) := To_stdlogicvector(X"00");
	mem(2031) := To_stdlogicvector(X"00");
	mem(2032) := To_stdlogicvector(X"00");
	mem(2033) := To_stdlogicvector(X"00");
	mem(2034) := To_stdlogicvector(X"00");
	mem(2035) := To_stdlogicvector(X"00");
	mem(2036) := To_stdlogicvector(X"00");
	mem(2037) := To_stdlogicvector(X"00");
	mem(2038) := To_stdlogicvector(X"00");
	mem(2039) := To_stdlogicvector(X"00");
	mem(2040) := To_stdlogicvector(X"00");
	mem(2041) := To_stdlogicvector(X"00");
	mem(2042) := To_stdlogicvector(X"00");
	mem(2043) := To_stdlogicvector(X"00");
	mem(2044) := To_stdlogicvector(X"00");
	mem(2045) := To_stdlogicvector(X"00");
	mem(2046) := To_stdlogicvector(X"00");
	mem(2047) := To_stdlogicvector(X"00");
	mem(2048) := To_stdlogicvector(X"00");
	mem(2049) := To_stdlogicvector(X"00");
	mem(2050) := To_stdlogicvector(X"00");
	mem(2051) := To_stdlogicvector(X"00");
	mem(2052) := To_stdlogicvector(X"00");
	mem(2053) := To_stdlogicvector(X"00");
	mem(2054) := To_stdlogicvector(X"00");
	mem(2055) := To_stdlogicvector(X"00");
	mem(2056) := To_stdlogicvector(X"00");
	mem(2057) := To_stdlogicvector(X"00");
	mem(2058) := To_stdlogicvector(X"00");
	mem(2059) := To_stdlogicvector(X"00");
	mem(2060) := To_stdlogicvector(X"00");
	mem(2061) := To_stdlogicvector(X"00");
	mem(2062) := To_stdlogicvector(X"00");
	mem(2063) := To_stdlogicvector(X"00");
	mem(2064) := To_stdlogicvector(X"00");
	mem(2065) := To_stdlogicvector(X"00");
	mem(2066) := To_stdlogicvector(X"00");
	mem(2067) := To_stdlogicvector(X"00");
	mem(2068) := To_stdlogicvector(X"00");
	mem(2069) := To_stdlogicvector(X"00");
	mem(2070) := To_stdlogicvector(X"00");
	mem(2071) := To_stdlogicvector(X"00");
	mem(2072) := To_stdlogicvector(X"00");
	mem(2073) := To_stdlogicvector(X"00");
	mem(2074) := To_stdlogicvector(X"00");
	mem(2075) := To_stdlogicvector(X"00");
	mem(2076) := To_stdlogicvector(X"00");
	mem(2077) := To_stdlogicvector(X"00");
	mem(2078) := To_stdlogicvector(X"00");
	mem(2079) := To_stdlogicvector(X"00");
	mem(2080) := To_stdlogicvector(X"00");
	mem(2081) := To_stdlogicvector(X"00");
	mem(2082) := To_stdlogicvector(X"00");
	mem(2083) := To_stdlogicvector(X"00");
	mem(2084) := To_stdlogicvector(X"00");
	mem(2085) := To_stdlogicvector(X"00");
	mem(2086) := To_stdlogicvector(X"00");
	mem(2087) := To_stdlogicvector(X"00");
	mem(2088) := To_stdlogicvector(X"00");
	mem(2089) := To_stdlogicvector(X"00");
	mem(2090) := To_stdlogicvector(X"00");
	mem(2091) := To_stdlogicvector(X"00");
	mem(2092) := To_stdlogicvector(X"00");
	mem(2093) := To_stdlogicvector(X"00");
	mem(2094) := To_stdlogicvector(X"00");
	mem(2095) := To_stdlogicvector(X"00");
	mem(2096) := To_stdlogicvector(X"00");
	mem(2097) := To_stdlogicvector(X"00");
	mem(2098) := To_stdlogicvector(X"00");
	mem(2099) := To_stdlogicvector(X"00");
	mem(2100) := To_stdlogicvector(X"00");
	mem(2101) := To_stdlogicvector(X"00");
	mem(2102) := To_stdlogicvector(X"00");
	mem(2103) := To_stdlogicvector(X"00");
	mem(2104) := To_stdlogicvector(X"00");
	mem(2105) := To_stdlogicvector(X"00");
	mem(2106) := To_stdlogicvector(X"00");
	mem(2107) := To_stdlogicvector(X"00");
	mem(2108) := To_stdlogicvector(X"00");
	mem(2109) := To_stdlogicvector(X"00");
	mem(2110) := To_stdlogicvector(X"00");
	mem(2111) := To_stdlogicvector(X"00");
	mem(2112) := To_stdlogicvector(X"00");
	mem(2113) := To_stdlogicvector(X"00");
	mem(2114) := To_stdlogicvector(X"00");
	mem(2115) := To_stdlogicvector(X"00");
	mem(2116) := To_stdlogicvector(X"00");
	mem(2117) := To_stdlogicvector(X"00");
	mem(2118) := To_stdlogicvector(X"00");
	mem(2119) := To_stdlogicvector(X"00");
	mem(2120) := To_stdlogicvector(X"00");
	mem(2121) := To_stdlogicvector(X"00");
	mem(2122) := To_stdlogicvector(X"00");
	mem(2123) := To_stdlogicvector(X"00");
	mem(2124) := To_stdlogicvector(X"00");
	mem(2125) := To_stdlogicvector(X"00");
	mem(2126) := To_stdlogicvector(X"00");
	mem(2127) := To_stdlogicvector(X"00");
	mem(2128) := To_stdlogicvector(X"00");
	mem(2129) := To_stdlogicvector(X"00");
	mem(2130) := To_stdlogicvector(X"00");
	mem(2131) := To_stdlogicvector(X"00");
	mem(2132) := To_stdlogicvector(X"00");
	mem(2133) := To_stdlogicvector(X"00");
	mem(2134) := To_stdlogicvector(X"00");
	mem(2135) := To_stdlogicvector(X"00");
	mem(2136) := To_stdlogicvector(X"00");
	mem(2137) := To_stdlogicvector(X"00");
	mem(2138) := To_stdlogicvector(X"00");
	mem(2139) := To_stdlogicvector(X"00");
	mem(2140) := To_stdlogicvector(X"00");
	mem(2141) := To_stdlogicvector(X"00");
	mem(2142) := To_stdlogicvector(X"00");
	mem(2143) := To_stdlogicvector(X"00");
	mem(2144) := To_stdlogicvector(X"00");
	mem(2145) := To_stdlogicvector(X"00");
	mem(2146) := To_stdlogicvector(X"00");
	mem(2147) := To_stdlogicvector(X"00");
	mem(2148) := To_stdlogicvector(X"00");
	mem(2149) := To_stdlogicvector(X"00");
	mem(2150) := To_stdlogicvector(X"00");
	mem(2151) := To_stdlogicvector(X"00");
	mem(2152) := To_stdlogicvector(X"00");
	mem(2153) := To_stdlogicvector(X"00");
	mem(2154) := To_stdlogicvector(X"00");
	mem(2155) := To_stdlogicvector(X"00");
	mem(2156) := To_stdlogicvector(X"00");
	mem(2157) := To_stdlogicvector(X"00");
	mem(2158) := To_stdlogicvector(X"00");
	mem(2159) := To_stdlogicvector(X"00");
	mem(2160) := To_stdlogicvector(X"00");
	mem(2161) := To_stdlogicvector(X"00");
	mem(2162) := To_stdlogicvector(X"00");
	mem(2163) := To_stdlogicvector(X"00");
	mem(2164) := To_stdlogicvector(X"00");
	mem(2165) := To_stdlogicvector(X"00");
	mem(2166) := To_stdlogicvector(X"00");
	mem(2167) := To_stdlogicvector(X"00");
	mem(2168) := To_stdlogicvector(X"00");
	mem(2169) := To_stdlogicvector(X"00");
	mem(2170) := To_stdlogicvector(X"00");
	mem(2171) := To_stdlogicvector(X"00");
	mem(2172) := To_stdlogicvector(X"00");
	mem(2173) := To_stdlogicvector(X"00");
	mem(2174) := To_stdlogicvector(X"00");
	mem(2175) := To_stdlogicvector(X"00");
	mem(2176) := To_stdlogicvector(X"00");
	mem(2177) := To_stdlogicvector(X"00");
	mem(2178) := To_stdlogicvector(X"00");
	mem(2179) := To_stdlogicvector(X"00");
	mem(2180) := To_stdlogicvector(X"00");
	mem(2181) := To_stdlogicvector(X"00");
	mem(2182) := To_stdlogicvector(X"00");
	mem(2183) := To_stdlogicvector(X"00");
	mem(2184) := To_stdlogicvector(X"00");
	mem(2185) := To_stdlogicvector(X"00");
	mem(2186) := To_stdlogicvector(X"00");
	mem(2187) := To_stdlogicvector(X"00");
	mem(2188) := To_stdlogicvector(X"00");
	mem(2189) := To_stdlogicvector(X"00");
	mem(2190) := To_stdlogicvector(X"00");
	mem(2191) := To_stdlogicvector(X"00");
	mem(2192) := To_stdlogicvector(X"00");
	mem(2193) := To_stdlogicvector(X"00");
	mem(2194) := To_stdlogicvector(X"00");
	mem(2195) := To_stdlogicvector(X"00");
	mem(2196) := To_stdlogicvector(X"00");
	mem(2197) := To_stdlogicvector(X"00");
	mem(2198) := To_stdlogicvector(X"00");
	mem(2199) := To_stdlogicvector(X"00");
	mem(2200) := To_stdlogicvector(X"00");
	mem(2201) := To_stdlogicvector(X"00");
	mem(2202) := To_stdlogicvector(X"00");
	mem(2203) := To_stdlogicvector(X"00");
	mem(2204) := To_stdlogicvector(X"00");
	mem(2205) := To_stdlogicvector(X"00");
	mem(2206) := To_stdlogicvector(X"00");
	mem(2207) := To_stdlogicvector(X"00");
	mem(2208) := To_stdlogicvector(X"00");
	mem(2209) := To_stdlogicvector(X"00");
	mem(2210) := To_stdlogicvector(X"00");
	mem(2211) := To_stdlogicvector(X"00");
	mem(2212) := To_stdlogicvector(X"00");
	mem(2213) := To_stdlogicvector(X"00");
	mem(2214) := To_stdlogicvector(X"00");
	mem(2215) := To_stdlogicvector(X"00");
	mem(2216) := To_stdlogicvector(X"00");
	mem(2217) := To_stdlogicvector(X"00");
	mem(2218) := To_stdlogicvector(X"00");
	mem(2219) := To_stdlogicvector(X"00");
	mem(2220) := To_stdlogicvector(X"00");
	mem(2221) := To_stdlogicvector(X"00");
	mem(2222) := To_stdlogicvector(X"00");
	mem(2223) := To_stdlogicvector(X"00");
	mem(2224) := To_stdlogicvector(X"00");
	mem(2225) := To_stdlogicvector(X"00");
	mem(2226) := To_stdlogicvector(X"00");
	mem(2227) := To_stdlogicvector(X"00");
	mem(2228) := To_stdlogicvector(X"00");
	mem(2229) := To_stdlogicvector(X"00");
	mem(2230) := To_stdlogicvector(X"00");
	mem(2231) := To_stdlogicvector(X"00");
	mem(2232) := To_stdlogicvector(X"00");
	mem(2233) := To_stdlogicvector(X"00");
	mem(2234) := To_stdlogicvector(X"00");
	mem(2235) := To_stdlogicvector(X"00");
	mem(2236) := To_stdlogicvector(X"00");
	mem(2237) := To_stdlogicvector(X"00");
	mem(2238) := To_stdlogicvector(X"00");
	mem(2239) := To_stdlogicvector(X"00");
	mem(2240) := To_stdlogicvector(X"00");
	mem(2241) := To_stdlogicvector(X"00");
	mem(2242) := To_stdlogicvector(X"00");
	mem(2243) := To_stdlogicvector(X"00");
	mem(2244) := To_stdlogicvector(X"00");
	mem(2245) := To_stdlogicvector(X"00");
	mem(2246) := To_stdlogicvector(X"00");
	mem(2247) := To_stdlogicvector(X"00");
	mem(2248) := To_stdlogicvector(X"00");
	mem(2249) := To_stdlogicvector(X"00");
	mem(2250) := To_stdlogicvector(X"00");
	mem(2251) := To_stdlogicvector(X"00");
	mem(2252) := To_stdlogicvector(X"00");
	mem(2253) := To_stdlogicvector(X"00");
	mem(2254) := To_stdlogicvector(X"00");
	mem(2255) := To_stdlogicvector(X"00");
	mem(2256) := To_stdlogicvector(X"00");
	mem(2257) := To_stdlogicvector(X"00");
	mem(2258) := To_stdlogicvector(X"00");
	mem(2259) := To_stdlogicvector(X"00");
	mem(2260) := To_stdlogicvector(X"00");
	mem(2261) := To_stdlogicvector(X"00");
	mem(2262) := To_stdlogicvector(X"00");
	mem(2263) := To_stdlogicvector(X"00");
	mem(2264) := To_stdlogicvector(X"00");
	mem(2265) := To_stdlogicvector(X"00");
	mem(2266) := To_stdlogicvector(X"00");
	mem(2267) := To_stdlogicvector(X"00");
	mem(2268) := To_stdlogicvector(X"00");
	mem(2269) := To_stdlogicvector(X"00");
	mem(2270) := To_stdlogicvector(X"00");
	mem(2271) := To_stdlogicvector(X"00");
	mem(2272) := To_stdlogicvector(X"00");
	mem(2273) := To_stdlogicvector(X"00");
	mem(2274) := To_stdlogicvector(X"00");
	mem(2275) := To_stdlogicvector(X"00");
	mem(2276) := To_stdlogicvector(X"00");
	mem(2277) := To_stdlogicvector(X"00");
	mem(2278) := To_stdlogicvector(X"00");
	mem(2279) := To_stdlogicvector(X"00");
	mem(2280) := To_stdlogicvector(X"00");
	mem(2281) := To_stdlogicvector(X"00");
	mem(2282) := To_stdlogicvector(X"00");
	mem(2283) := To_stdlogicvector(X"00");
	mem(2284) := To_stdlogicvector(X"00");
	mem(2285) := To_stdlogicvector(X"00");
	mem(2286) := To_stdlogicvector(X"00");
	mem(2287) := To_stdlogicvector(X"00");
	mem(2288) := To_stdlogicvector(X"00");
	mem(2289) := To_stdlogicvector(X"00");
	mem(2290) := To_stdlogicvector(X"00");
	mem(2291) := To_stdlogicvector(X"00");
	mem(2292) := To_stdlogicvector(X"00");
	mem(2293) := To_stdlogicvector(X"00");
	mem(2294) := To_stdlogicvector(X"00");
	mem(2295) := To_stdlogicvector(X"00");
	mem(2296) := To_stdlogicvector(X"00");
	mem(2297) := To_stdlogicvector(X"00");
	mem(2298) := To_stdlogicvector(X"00");
	mem(2299) := To_stdlogicvector(X"00");
	mem(2300) := To_stdlogicvector(X"00");
	mem(2301) := To_stdlogicvector(X"00");
	mem(2302) := To_stdlogicvector(X"00");
	mem(2303) := To_stdlogicvector(X"00");
	mem(2304) := To_stdlogicvector(X"00");
	mem(2305) := To_stdlogicvector(X"00");
	mem(2306) := To_stdlogicvector(X"00");
	mem(2307) := To_stdlogicvector(X"00");
	mem(2308) := To_stdlogicvector(X"00");
	mem(2309) := To_stdlogicvector(X"00");
	mem(2310) := To_stdlogicvector(X"00");
	mem(2311) := To_stdlogicvector(X"00");
	mem(2312) := To_stdlogicvector(X"00");
	mem(2313) := To_stdlogicvector(X"00");
	mem(2314) := To_stdlogicvector(X"00");
	mem(2315) := To_stdlogicvector(X"00");
	mem(2316) := To_stdlogicvector(X"00");
	mem(2317) := To_stdlogicvector(X"00");
	mem(2318) := To_stdlogicvector(X"00");
	mem(2319) := To_stdlogicvector(X"00");
	mem(2320) := To_stdlogicvector(X"00");
	mem(2321) := To_stdlogicvector(X"00");
	mem(2322) := To_stdlogicvector(X"00");
	mem(2323) := To_stdlogicvector(X"00");
	mem(2324) := To_stdlogicvector(X"00");
	mem(2325) := To_stdlogicvector(X"00");
	mem(2326) := To_stdlogicvector(X"00");
	mem(2327) := To_stdlogicvector(X"00");
	mem(2328) := To_stdlogicvector(X"00");
	mem(2329) := To_stdlogicvector(X"00");
	mem(2330) := To_stdlogicvector(X"00");
	mem(2331) := To_stdlogicvector(X"00");
	mem(2332) := To_stdlogicvector(X"00");
	mem(2333) := To_stdlogicvector(X"00");
	mem(2334) := To_stdlogicvector(X"00");
	mem(2335) := To_stdlogicvector(X"00");
	mem(2336) := To_stdlogicvector(X"00");
	mem(2337) := To_stdlogicvector(X"00");
	mem(2338) := To_stdlogicvector(X"00");
	mem(2339) := To_stdlogicvector(X"00");
	mem(2340) := To_stdlogicvector(X"00");
	mem(2341) := To_stdlogicvector(X"00");
	mem(2342) := To_stdlogicvector(X"00");
	mem(2343) := To_stdlogicvector(X"00");
	mem(2344) := To_stdlogicvector(X"00");
	mem(2345) := To_stdlogicvector(X"00");
	mem(2346) := To_stdlogicvector(X"00");
	mem(2347) := To_stdlogicvector(X"00");
	mem(2348) := To_stdlogicvector(X"00");
	mem(2349) := To_stdlogicvector(X"00");
	mem(2350) := To_stdlogicvector(X"00");
	mem(2351) := To_stdlogicvector(X"00");
	mem(2352) := To_stdlogicvector(X"00");
	mem(2353) := To_stdlogicvector(X"00");
	mem(2354) := To_stdlogicvector(X"00");
	mem(2355) := To_stdlogicvector(X"00");
	mem(2356) := To_stdlogicvector(X"00");
	mem(2357) := To_stdlogicvector(X"00");
	mem(2358) := To_stdlogicvector(X"00");
	mem(2359) := To_stdlogicvector(X"00");
	mem(2360) := To_stdlogicvector(X"00");
	mem(2361) := To_stdlogicvector(X"00");
	mem(2362) := To_stdlogicvector(X"00");
	mem(2363) := To_stdlogicvector(X"00");
	mem(2364) := To_stdlogicvector(X"00");
	mem(2365) := To_stdlogicvector(X"00");
	mem(2366) := To_stdlogicvector(X"00");
	mem(2367) := To_stdlogicvector(X"00");
	mem(2368) := To_stdlogicvector(X"00");
	mem(2369) := To_stdlogicvector(X"00");
	mem(2370) := To_stdlogicvector(X"00");
	mem(2371) := To_stdlogicvector(X"00");
	mem(2372) := To_stdlogicvector(X"00");
	mem(2373) := To_stdlogicvector(X"00");
	mem(2374) := To_stdlogicvector(X"00");
	mem(2375) := To_stdlogicvector(X"00");
	mem(2376) := To_stdlogicvector(X"00");
	mem(2377) := To_stdlogicvector(X"00");
	mem(2378) := To_stdlogicvector(X"00");
	mem(2379) := To_stdlogicvector(X"00");
	mem(2380) := To_stdlogicvector(X"00");
	mem(2381) := To_stdlogicvector(X"00");
	mem(2382) := To_stdlogicvector(X"00");
	mem(2383) := To_stdlogicvector(X"00");
	mem(2384) := To_stdlogicvector(X"00");
	mem(2385) := To_stdlogicvector(X"00");
	mem(2386) := To_stdlogicvector(X"00");
	mem(2387) := To_stdlogicvector(X"00");
	mem(2388) := To_stdlogicvector(X"00");
	mem(2389) := To_stdlogicvector(X"00");
	mem(2390) := To_stdlogicvector(X"00");
	mem(2391) := To_stdlogicvector(X"00");
	mem(2392) := To_stdlogicvector(X"00");
	mem(2393) := To_stdlogicvector(X"00");
	mem(2394) := To_stdlogicvector(X"00");
	mem(2395) := To_stdlogicvector(X"00");
	mem(2396) := To_stdlogicvector(X"00");
	mem(2397) := To_stdlogicvector(X"00");
	mem(2398) := To_stdlogicvector(X"00");
	mem(2399) := To_stdlogicvector(X"00");
	mem(2400) := To_stdlogicvector(X"00");
	mem(2401) := To_stdlogicvector(X"00");
	mem(2402) := To_stdlogicvector(X"00");
	mem(2403) := To_stdlogicvector(X"00");
	mem(2404) := To_stdlogicvector(X"00");
	mem(2405) := To_stdlogicvector(X"00");
	mem(2406) := To_stdlogicvector(X"00");
	mem(2407) := To_stdlogicvector(X"00");
	mem(2408) := To_stdlogicvector(X"00");
	mem(2409) := To_stdlogicvector(X"00");
	mem(2410) := To_stdlogicvector(X"00");
	mem(2411) := To_stdlogicvector(X"00");
	mem(2412) := To_stdlogicvector(X"00");
	mem(2413) := To_stdlogicvector(X"00");
	mem(2414) := To_stdlogicvector(X"00");
	mem(2415) := To_stdlogicvector(X"00");
	mem(2416) := To_stdlogicvector(X"00");
	mem(2417) := To_stdlogicvector(X"00");
	mem(2418) := To_stdlogicvector(X"00");
	mem(2419) := To_stdlogicvector(X"00");
	mem(2420) := To_stdlogicvector(X"00");
	mem(2421) := To_stdlogicvector(X"00");
	mem(2422) := To_stdlogicvector(X"00");
	mem(2423) := To_stdlogicvector(X"00");
	mem(2424) := To_stdlogicvector(X"00");
	mem(2425) := To_stdlogicvector(X"00");
	mem(2426) := To_stdlogicvector(X"00");
	mem(2427) := To_stdlogicvector(X"00");
	mem(2428) := To_stdlogicvector(X"00");
	mem(2429) := To_stdlogicvector(X"00");
	mem(2430) := To_stdlogicvector(X"00");
	mem(2431) := To_stdlogicvector(X"00");
	mem(2432) := To_stdlogicvector(X"00");
	mem(2433) := To_stdlogicvector(X"00");
	mem(2434) := To_stdlogicvector(X"00");
	mem(2435) := To_stdlogicvector(X"00");
	mem(2436) := To_stdlogicvector(X"00");
	mem(2437) := To_stdlogicvector(X"00");
	mem(2438) := To_stdlogicvector(X"00");
	mem(2439) := To_stdlogicvector(X"00");
	mem(2440) := To_stdlogicvector(X"00");
	mem(2441) := To_stdlogicvector(X"00");
	mem(2442) := To_stdlogicvector(X"00");
	mem(2443) := To_stdlogicvector(X"00");
	mem(2444) := To_stdlogicvector(X"00");
	mem(2445) := To_stdlogicvector(X"00");
	mem(2446) := To_stdlogicvector(X"00");
	mem(2447) := To_stdlogicvector(X"00");
	mem(2448) := To_stdlogicvector(X"00");
	mem(2449) := To_stdlogicvector(X"00");
	mem(2450) := To_stdlogicvector(X"00");
	mem(2451) := To_stdlogicvector(X"00");
	mem(2452) := To_stdlogicvector(X"00");
	mem(2453) := To_stdlogicvector(X"00");
	mem(2454) := To_stdlogicvector(X"00");
	mem(2455) := To_stdlogicvector(X"00");
	mem(2456) := To_stdlogicvector(X"00");
	mem(2457) := To_stdlogicvector(X"00");
	mem(2458) := To_stdlogicvector(X"00");
	mem(2459) := To_stdlogicvector(X"00");
	mem(2460) := To_stdlogicvector(X"00");
	mem(2461) := To_stdlogicvector(X"00");
	mem(2462) := To_stdlogicvector(X"00");
	mem(2463) := To_stdlogicvector(X"00");
	mem(2464) := To_stdlogicvector(X"00");
	mem(2465) := To_stdlogicvector(X"00");
	mem(2466) := To_stdlogicvector(X"00");
	mem(2467) := To_stdlogicvector(X"00");
	mem(2468) := To_stdlogicvector(X"00");
	mem(2469) := To_stdlogicvector(X"00");
	mem(2470) := To_stdlogicvector(X"00");
	mem(2471) := To_stdlogicvector(X"00");
	mem(2472) := To_stdlogicvector(X"00");
	mem(2473) := To_stdlogicvector(X"00");
	mem(2474) := To_stdlogicvector(X"00");
	mem(2475) := To_stdlogicvector(X"00");
	mem(2476) := To_stdlogicvector(X"00");
	mem(2477) := To_stdlogicvector(X"00");
	mem(2478) := To_stdlogicvector(X"00");
	mem(2479) := To_stdlogicvector(X"00");
	mem(2480) := To_stdlogicvector(X"00");
	mem(2481) := To_stdlogicvector(X"00");
	mem(2482) := To_stdlogicvector(X"00");
	mem(2483) := To_stdlogicvector(X"00");
	mem(2484) := To_stdlogicvector(X"00");
	mem(2485) := To_stdlogicvector(X"00");
	mem(2486) := To_stdlogicvector(X"00");
	mem(2487) := To_stdlogicvector(X"00");
	mem(2488) := To_stdlogicvector(X"00");
	mem(2489) := To_stdlogicvector(X"00");
	mem(2490) := To_stdlogicvector(X"00");
	mem(2491) := To_stdlogicvector(X"00");
	mem(2492) := To_stdlogicvector(X"00");
	mem(2493) := To_stdlogicvector(X"00");
	mem(2494) := To_stdlogicvector(X"00");
	mem(2495) := To_stdlogicvector(X"00");
	mem(2496) := To_stdlogicvector(X"00");
	mem(2497) := To_stdlogicvector(X"00");
	mem(2498) := To_stdlogicvector(X"00");
	mem(2499) := To_stdlogicvector(X"00");
	mem(2500) := To_stdlogicvector(X"00");
	mem(2501) := To_stdlogicvector(X"00");
	mem(2502) := To_stdlogicvector(X"00");
	mem(2503) := To_stdlogicvector(X"00");
	mem(2504) := To_stdlogicvector(X"00");
	mem(2505) := To_stdlogicvector(X"00");
	mem(2506) := To_stdlogicvector(X"00");
	mem(2507) := To_stdlogicvector(X"00");
	mem(2508) := To_stdlogicvector(X"00");
	mem(2509) := To_stdlogicvector(X"00");
	mem(2510) := To_stdlogicvector(X"00");
	mem(2511) := To_stdlogicvector(X"00");
	mem(2512) := To_stdlogicvector(X"00");
	mem(2513) := To_stdlogicvector(X"00");
	mem(2514) := To_stdlogicvector(X"00");
	mem(2515) := To_stdlogicvector(X"00");
	mem(2516) := To_stdlogicvector(X"00");
	mem(2517) := To_stdlogicvector(X"00");
	mem(2518) := To_stdlogicvector(X"00");
	mem(2519) := To_stdlogicvector(X"00");
	mem(2520) := To_stdlogicvector(X"00");
	mem(2521) := To_stdlogicvector(X"00");
	mem(2522) := To_stdlogicvector(X"00");
	mem(2523) := To_stdlogicvector(X"00");
	mem(2524) := To_stdlogicvector(X"00");
	mem(2525) := To_stdlogicvector(X"00");
	mem(2526) := To_stdlogicvector(X"00");
	mem(2527) := To_stdlogicvector(X"00");
	mem(2528) := To_stdlogicvector(X"00");
	mem(2529) := To_stdlogicvector(X"00");
	mem(2530) := To_stdlogicvector(X"00");
	mem(2531) := To_stdlogicvector(X"00");
	mem(2532) := To_stdlogicvector(X"00");
	mem(2533) := To_stdlogicvector(X"00");
	mem(2534) := To_stdlogicvector(X"00");
	mem(2535) := To_stdlogicvector(X"00");
	mem(2536) := To_stdlogicvector(X"00");
	mem(2537) := To_stdlogicvector(X"00");
	mem(2538) := To_stdlogicvector(X"00");
	mem(2539) := To_stdlogicvector(X"00");
	mem(2540) := To_stdlogicvector(X"00");
	mem(2541) := To_stdlogicvector(X"00");
	mem(2542) := To_stdlogicvector(X"00");
	mem(2543) := To_stdlogicvector(X"00");
	mem(2544) := To_stdlogicvector(X"00");
	mem(2545) := To_stdlogicvector(X"00");
	mem(2546) := To_stdlogicvector(X"00");
	mem(2547) := To_stdlogicvector(X"00");
	mem(2548) := To_stdlogicvector(X"00");
	mem(2549) := To_stdlogicvector(X"00");
	mem(2550) := To_stdlogicvector(X"00");
	mem(2551) := To_stdlogicvector(X"00");
	mem(2552) := To_stdlogicvector(X"00");
	mem(2553) := To_stdlogicvector(X"00");
	mem(2554) := To_stdlogicvector(X"00");
	mem(2555) := To_stdlogicvector(X"00");
	mem(2556) := To_stdlogicvector(X"00");
	mem(2557) := To_stdlogicvector(X"00");
	mem(2558) := To_stdlogicvector(X"00");
	mem(2559) := To_stdlogicvector(X"00");
	mem(2560) := To_stdlogicvector(X"00");
	mem(2561) := To_stdlogicvector(X"00");
	mem(2562) := To_stdlogicvector(X"00");
	mem(2563) := To_stdlogicvector(X"00");
	mem(2564) := To_stdlogicvector(X"00");
	mem(2565) := To_stdlogicvector(X"00");
	mem(2566) := To_stdlogicvector(X"00");
	mem(2567) := To_stdlogicvector(X"00");
	mem(2568) := To_stdlogicvector(X"00");
	mem(2569) := To_stdlogicvector(X"00");
	mem(2570) := To_stdlogicvector(X"00");
	mem(2571) := To_stdlogicvector(X"00");
	mem(2572) := To_stdlogicvector(X"00");
	mem(2573) := To_stdlogicvector(X"00");
	mem(2574) := To_stdlogicvector(X"00");
	mem(2575) := To_stdlogicvector(X"00");
	mem(2576) := To_stdlogicvector(X"00");
	mem(2577) := To_stdlogicvector(X"00");
	mem(2578) := To_stdlogicvector(X"00");
	mem(2579) := To_stdlogicvector(X"00");
	mem(2580) := To_stdlogicvector(X"00");
	mem(2581) := To_stdlogicvector(X"00");
	mem(2582) := To_stdlogicvector(X"00");
	mem(2583) := To_stdlogicvector(X"00");
	mem(2584) := To_stdlogicvector(X"00");
	mem(2585) := To_stdlogicvector(X"00");
	mem(2586) := To_stdlogicvector(X"00");
	mem(2587) := To_stdlogicvector(X"00");
	mem(2588) := To_stdlogicvector(X"00");
	mem(2589) := To_stdlogicvector(X"00");
	mem(2590) := To_stdlogicvector(X"00");
	mem(2591) := To_stdlogicvector(X"00");
	mem(2592) := To_stdlogicvector(X"00");
	mem(2593) := To_stdlogicvector(X"00");
	mem(2594) := To_stdlogicvector(X"00");
	mem(2595) := To_stdlogicvector(X"00");
	mem(2596) := To_stdlogicvector(X"00");
	mem(2597) := To_stdlogicvector(X"00");
	mem(2598) := To_stdlogicvector(X"00");
	mem(2599) := To_stdlogicvector(X"00");
	mem(2600) := To_stdlogicvector(X"00");
	mem(2601) := To_stdlogicvector(X"00");
	mem(2602) := To_stdlogicvector(X"00");
	mem(2603) := To_stdlogicvector(X"00");
	mem(2604) := To_stdlogicvector(X"00");
	mem(2605) := To_stdlogicvector(X"00");
	mem(2606) := To_stdlogicvector(X"00");
	mem(2607) := To_stdlogicvector(X"00");
	mem(2608) := To_stdlogicvector(X"00");
	mem(2609) := To_stdlogicvector(X"00");
	mem(2610) := To_stdlogicvector(X"00");
	mem(2611) := To_stdlogicvector(X"00");
	mem(2612) := To_stdlogicvector(X"00");
	mem(2613) := To_stdlogicvector(X"00");
	mem(2614) := To_stdlogicvector(X"00");
	mem(2615) := To_stdlogicvector(X"00");
	mem(2616) := To_stdlogicvector(X"00");
	mem(2617) := To_stdlogicvector(X"00");
	mem(2618) := To_stdlogicvector(X"00");
	mem(2619) := To_stdlogicvector(X"00");
	mem(2620) := To_stdlogicvector(X"00");
	mem(2621) := To_stdlogicvector(X"00");
	mem(2622) := To_stdlogicvector(X"00");
	mem(2623) := To_stdlogicvector(X"00");
	mem(2624) := To_stdlogicvector(X"00");
	mem(2625) := To_stdlogicvector(X"00");
	mem(2626) := To_stdlogicvector(X"00");
	mem(2627) := To_stdlogicvector(X"00");
	mem(2628) := To_stdlogicvector(X"00");
	mem(2629) := To_stdlogicvector(X"00");
	mem(2630) := To_stdlogicvector(X"00");
	mem(2631) := To_stdlogicvector(X"00");
	mem(2632) := To_stdlogicvector(X"00");
	mem(2633) := To_stdlogicvector(X"00");
	mem(2634) := To_stdlogicvector(X"00");
	mem(2635) := To_stdlogicvector(X"00");
	mem(2636) := To_stdlogicvector(X"00");
	mem(2637) := To_stdlogicvector(X"00");
	mem(2638) := To_stdlogicvector(X"00");
	mem(2639) := To_stdlogicvector(X"00");
	mem(2640) := To_stdlogicvector(X"00");
	mem(2641) := To_stdlogicvector(X"00");
	mem(2642) := To_stdlogicvector(X"00");
	mem(2643) := To_stdlogicvector(X"00");
	mem(2644) := To_stdlogicvector(X"00");
	mem(2645) := To_stdlogicvector(X"00");
	mem(2646) := To_stdlogicvector(X"00");
	mem(2647) := To_stdlogicvector(X"00");
	mem(2648) := To_stdlogicvector(X"00");
	mem(2649) := To_stdlogicvector(X"00");
	mem(2650) := To_stdlogicvector(X"00");
	mem(2651) := To_stdlogicvector(X"00");
	mem(2652) := To_stdlogicvector(X"00");
	mem(2653) := To_stdlogicvector(X"00");
	mem(2654) := To_stdlogicvector(X"00");
	mem(2655) := To_stdlogicvector(X"00");
	mem(2656) := To_stdlogicvector(X"00");
	mem(2657) := To_stdlogicvector(X"00");
	mem(2658) := To_stdlogicvector(X"00");
	mem(2659) := To_stdlogicvector(X"00");
	mem(2660) := To_stdlogicvector(X"00");
	mem(2661) := To_stdlogicvector(X"00");
	mem(2662) := To_stdlogicvector(X"00");
	mem(2663) := To_stdlogicvector(X"00");
	mem(2664) := To_stdlogicvector(X"00");
	mem(2665) := To_stdlogicvector(X"00");
	mem(2666) := To_stdlogicvector(X"00");
	mem(2667) := To_stdlogicvector(X"00");
	mem(2668) := To_stdlogicvector(X"00");
	mem(2669) := To_stdlogicvector(X"00");
	mem(2670) := To_stdlogicvector(X"00");
	mem(2671) := To_stdlogicvector(X"00");
	mem(2672) := To_stdlogicvector(X"00");
	mem(2673) := To_stdlogicvector(X"00");
	mem(2674) := To_stdlogicvector(X"00");
	mem(2675) := To_stdlogicvector(X"00");
	mem(2676) := To_stdlogicvector(X"00");
	mem(2677) := To_stdlogicvector(X"00");
	mem(2678) := To_stdlogicvector(X"00");
	mem(2679) := To_stdlogicvector(X"00");
	mem(2680) := To_stdlogicvector(X"00");
	mem(2681) := To_stdlogicvector(X"00");
	mem(2682) := To_stdlogicvector(X"00");
	mem(2683) := To_stdlogicvector(X"00");
	mem(2684) := To_stdlogicvector(X"00");
	mem(2685) := To_stdlogicvector(X"00");
	mem(2686) := To_stdlogicvector(X"00");
	mem(2687) := To_stdlogicvector(X"00");
	mem(2688) := To_stdlogicvector(X"00");
	mem(2689) := To_stdlogicvector(X"00");
	mem(2690) := To_stdlogicvector(X"00");
	mem(2691) := To_stdlogicvector(X"00");
	mem(2692) := To_stdlogicvector(X"00");
	mem(2693) := To_stdlogicvector(X"00");
	mem(2694) := To_stdlogicvector(X"00");
	mem(2695) := To_stdlogicvector(X"00");
	mem(2696) := To_stdlogicvector(X"00");
	mem(2697) := To_stdlogicvector(X"00");
	mem(2698) := To_stdlogicvector(X"00");
	mem(2699) := To_stdlogicvector(X"00");
	mem(2700) := To_stdlogicvector(X"00");
	mem(2701) := To_stdlogicvector(X"00");
	mem(2702) := To_stdlogicvector(X"00");
	mem(2703) := To_stdlogicvector(X"00");
	mem(2704) := To_stdlogicvector(X"00");
	mem(2705) := To_stdlogicvector(X"00");
	mem(2706) := To_stdlogicvector(X"00");
	mem(2707) := To_stdlogicvector(X"00");
	mem(2708) := To_stdlogicvector(X"00");
	mem(2709) := To_stdlogicvector(X"00");
	mem(2710) := To_stdlogicvector(X"00");
	mem(2711) := To_stdlogicvector(X"00");
	mem(2712) := To_stdlogicvector(X"00");
	mem(2713) := To_stdlogicvector(X"00");
	mem(2714) := To_stdlogicvector(X"00");
	mem(2715) := To_stdlogicvector(X"00");
	mem(2716) := To_stdlogicvector(X"00");
	mem(2717) := To_stdlogicvector(X"00");
	mem(2718) := To_stdlogicvector(X"00");
	mem(2719) := To_stdlogicvector(X"00");
	mem(2720) := To_stdlogicvector(X"00");
	mem(2721) := To_stdlogicvector(X"00");
	mem(2722) := To_stdlogicvector(X"00");
	mem(2723) := To_stdlogicvector(X"00");
	mem(2724) := To_stdlogicvector(X"00");
	mem(2725) := To_stdlogicvector(X"00");
	mem(2726) := To_stdlogicvector(X"00");
	mem(2727) := To_stdlogicvector(X"00");
	mem(2728) := To_stdlogicvector(X"00");
	mem(2729) := To_stdlogicvector(X"00");
	mem(2730) := To_stdlogicvector(X"00");
	mem(2731) := To_stdlogicvector(X"00");
	mem(2732) := To_stdlogicvector(X"00");
	mem(2733) := To_stdlogicvector(X"00");
	mem(2734) := To_stdlogicvector(X"00");
	mem(2735) := To_stdlogicvector(X"00");
	mem(2736) := To_stdlogicvector(X"00");
	mem(2737) := To_stdlogicvector(X"00");
	mem(2738) := To_stdlogicvector(X"00");
	mem(2739) := To_stdlogicvector(X"00");
	mem(2740) := To_stdlogicvector(X"00");
	mem(2741) := To_stdlogicvector(X"00");
	mem(2742) := To_stdlogicvector(X"00");
	mem(2743) := To_stdlogicvector(X"00");
	mem(2744) := To_stdlogicvector(X"00");
	mem(2745) := To_stdlogicvector(X"00");
	mem(2746) := To_stdlogicvector(X"00");
	mem(2747) := To_stdlogicvector(X"00");
	mem(2748) := To_stdlogicvector(X"00");
	mem(2749) := To_stdlogicvector(X"00");
	mem(2750) := To_stdlogicvector(X"00");
	mem(2751) := To_stdlogicvector(X"00");
	mem(2752) := To_stdlogicvector(X"00");
	mem(2753) := To_stdlogicvector(X"00");
	mem(2754) := To_stdlogicvector(X"00");
	mem(2755) := To_stdlogicvector(X"00");
	mem(2756) := To_stdlogicvector(X"00");
	mem(2757) := To_stdlogicvector(X"00");
	mem(2758) := To_stdlogicvector(X"00");
	mem(2759) := To_stdlogicvector(X"00");
	mem(2760) := To_stdlogicvector(X"00");
	mem(2761) := To_stdlogicvector(X"00");
	mem(2762) := To_stdlogicvector(X"00");
	mem(2763) := To_stdlogicvector(X"00");
	mem(2764) := To_stdlogicvector(X"00");
	mem(2765) := To_stdlogicvector(X"00");
	mem(2766) := To_stdlogicvector(X"00");
	mem(2767) := To_stdlogicvector(X"00");
	mem(2768) := To_stdlogicvector(X"00");
	mem(2769) := To_stdlogicvector(X"00");
	mem(2770) := To_stdlogicvector(X"00");
	mem(2771) := To_stdlogicvector(X"00");
	mem(2772) := To_stdlogicvector(X"00");
	mem(2773) := To_stdlogicvector(X"00");
	mem(2774) := To_stdlogicvector(X"00");
	mem(2775) := To_stdlogicvector(X"00");
	mem(2776) := To_stdlogicvector(X"00");
	mem(2777) := To_stdlogicvector(X"00");
	mem(2778) := To_stdlogicvector(X"00");
	mem(2779) := To_stdlogicvector(X"00");
	mem(2780) := To_stdlogicvector(X"00");
	mem(2781) := To_stdlogicvector(X"00");
	mem(2782) := To_stdlogicvector(X"00");
	mem(2783) := To_stdlogicvector(X"00");
	mem(2784) := To_stdlogicvector(X"00");
	mem(2785) := To_stdlogicvector(X"00");
	mem(2786) := To_stdlogicvector(X"00");
	mem(2787) := To_stdlogicvector(X"00");
