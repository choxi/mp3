	mem(0) := To_stdlogicvector(X"07");
	mem(1) := To_stdlogicvector(X"E0");
	mem(2) := To_stdlogicvector(X"00");
	mem(3) := To_stdlogicvector(X"00");
	mem(4) := To_stdlogicvector(X"00");
	mem(5) := To_stdlogicvector(X"00");
	mem(6) := To_stdlogicvector(X"00");
	mem(7) := To_stdlogicvector(X"00");
	mem(8) := To_stdlogicvector(X"00");
	mem(9) := To_stdlogicvector(X"00");
	mem(10) := To_stdlogicvector(X"00");
	mem(11) := To_stdlogicvector(X"00");
	mem(12) := To_stdlogicvector(X"00");
	mem(13) := To_stdlogicvector(X"00");
	mem(14) := To_stdlogicvector(X"20");
	mem(15) := To_stdlogicvector(X"0E");
	mem(16) := To_stdlogicvector(X"00");
	mem(17) := To_stdlogicvector(X"00");
	mem(18) := To_stdlogicvector(X"70");
	mem(19) := To_stdlogicvector(X"00");
	mem(20) := To_stdlogicvector(X"0A");
	mem(21) := To_stdlogicvector(X"00");
	mem(22) := To_stdlogicvector(X"0F");
	mem(23) := To_stdlogicvector(X"27");
	mem(24) := To_stdlogicvector(X"2A");
	mem(25) := To_stdlogicvector(X"00");
	mem(26) := To_stdlogicvector(X"C8");
	mem(27) := To_stdlogicvector(X"BA");
	mem(28) := To_stdlogicvector(X"07");
	mem(29) := To_stdlogicvector(X"00");
	mem(30) := To_stdlogicvector(X"03");
	mem(31) := To_stdlogicvector(X"00");
	mem(32) := To_stdlogicvector(X"AD");
	mem(33) := To_stdlogicvector(X"0B");
	mem(34) := To_stdlogicvector(X"0D");
	mem(35) := To_stdlogicvector(X"0D");
	mem(36) := To_stdlogicvector(X"84");
	mem(37) := To_stdlogicvector(X"98");
	mem(38) := To_stdlogicvector(X"85");
	mem(39) := To_stdlogicvector(X"AE");
	mem(40) := To_stdlogicvector(X"60");
	mem(41) := To_stdlogicvector(X"54");
	mem(42) := To_stdlogicvector(X"05");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"46");
	mem(45) := To_stdlogicvector(X"06");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"00");
	mem(49) := To_stdlogicvector(X"00");
	mem(50) := To_stdlogicvector(X"00");
	mem(51) := To_stdlogicvector(X"00");
	mem(52) := To_stdlogicvector(X"00");
	mem(53) := To_stdlogicvector(X"00");
	mem(54) := To_stdlogicvector(X"00");
	mem(55) := To_stdlogicvector(X"00");
	mem(56) := To_stdlogicvector(X"00");
	mem(57) := To_stdlogicvector(X"00");
	mem(58) := To_stdlogicvector(X"00");
	mem(59) := To_stdlogicvector(X"00");
	mem(60) := To_stdlogicvector(X"00");
	mem(61) := To_stdlogicvector(X"00");
	mem(62) := To_stdlogicvector(X"00");
	mem(63) := To_stdlogicvector(X"00");
	mem(64) := To_stdlogicvector(X"00");
	mem(65) := To_stdlogicvector(X"00");
	mem(66) := To_stdlogicvector(X"00");
	mem(67) := To_stdlogicvector(X"00");
	mem(68) := To_stdlogicvector(X"00");
	mem(69) := To_stdlogicvector(X"00");
	mem(70) := To_stdlogicvector(X"00");
	mem(71) := To_stdlogicvector(X"00");
	mem(72) := To_stdlogicvector(X"00");
	mem(73) := To_stdlogicvector(X"00");
	mem(74) := To_stdlogicvector(X"00");
	mem(75) := To_stdlogicvector(X"00");
	mem(76) := To_stdlogicvector(X"00");
	mem(77) := To_stdlogicvector(X"00");
	mem(78) := To_stdlogicvector(X"1E");
	mem(79) := To_stdlogicvector(X"04");
	mem(80) := To_stdlogicvector(X"00");
	mem(81) := To_stdlogicvector(X"62");
	mem(82) := To_stdlogicvector(X"00");
	mem(83) := To_stdlogicvector(X"00");
	mem(84) := To_stdlogicvector(X"00");
	mem(85) := To_stdlogicvector(X"00");
	mem(86) := To_stdlogicvector(X"00");
	mem(87) := To_stdlogicvector(X"00");
	mem(88) := To_stdlogicvector(X"00");
	mem(89) := To_stdlogicvector(X"00");
	mem(90) := To_stdlogicvector(X"00");
	mem(91) := To_stdlogicvector(X"00");
	mem(92) := To_stdlogicvector(X"00");
	mem(93) := To_stdlogicvector(X"00");
	mem(94) := To_stdlogicvector(X"01");
	mem(95) := To_stdlogicvector(X"64");
	mem(96) := To_stdlogicvector(X"00");
	mem(97) := To_stdlogicvector(X"00");
	mem(98) := To_stdlogicvector(X"00");
	mem(99) := To_stdlogicvector(X"00");
	mem(100) := To_stdlogicvector(X"00");
	mem(101) := To_stdlogicvector(X"00");
	mem(102) := To_stdlogicvector(X"00");
	mem(103) := To_stdlogicvector(X"00");
	mem(104) := To_stdlogicvector(X"00");
	mem(105) := To_stdlogicvector(X"00");
	mem(106) := To_stdlogicvector(X"00");
	mem(107) := To_stdlogicvector(X"00");
	mem(108) := To_stdlogicvector(X"02");
	mem(109) := To_stdlogicvector(X"6E");
	mem(110) := To_stdlogicvector(X"00");
	mem(111) := To_stdlogicvector(X"00");
	mem(112) := To_stdlogicvector(X"00");
	mem(113) := To_stdlogicvector(X"00");
	mem(114) := To_stdlogicvector(X"00");
	mem(115) := To_stdlogicvector(X"00");
	mem(116) := To_stdlogicvector(X"00");
	mem(117) := To_stdlogicvector(X"00");
	mem(118) := To_stdlogicvector(X"00");
	mem(119) := To_stdlogicvector(X"00");
	mem(120) := To_stdlogicvector(X"00");
	mem(121) := To_stdlogicvector(X"00");
	mem(122) := To_stdlogicvector(X"87");
	mem(123) := To_stdlogicvector(X"12");
	mem(124) := To_stdlogicvector(X"00");
	mem(125) := To_stdlogicvector(X"00");
	mem(126) := To_stdlogicvector(X"00");
	mem(127) := To_stdlogicvector(X"00");
	mem(128) := To_stdlogicvector(X"00");
	mem(129) := To_stdlogicvector(X"00");
	mem(130) := To_stdlogicvector(X"00");
	mem(131) := To_stdlogicvector(X"00");
	mem(132) := To_stdlogicvector(X"00");
	mem(133) := To_stdlogicvector(X"00");
	mem(134) := To_stdlogicvector(X"00");
	mem(135) := To_stdlogicvector(X"00");
	mem(136) := To_stdlogicvector(X"7C");
	mem(137) := To_stdlogicvector(X"16");
	mem(138) := To_stdlogicvector(X"00");
	mem(139) := To_stdlogicvector(X"00");
	mem(140) := To_stdlogicvector(X"00");
	mem(141) := To_stdlogicvector(X"00");
	mem(142) := To_stdlogicvector(X"00");
	mem(143) := To_stdlogicvector(X"00");
	mem(144) := To_stdlogicvector(X"00");
	mem(145) := To_stdlogicvector(X"00");
	mem(146) := To_stdlogicvector(X"00");
	mem(147) := To_stdlogicvector(X"00");
	mem(148) := To_stdlogicvector(X"00");
	mem(149) := To_stdlogicvector(X"00");
	mem(150) := To_stdlogicvector(X"43");
	mem(151) := To_stdlogicvector(X"12");
	mem(152) := To_stdlogicvector(X"00");
	mem(153) := To_stdlogicvector(X"00");
	mem(154) := To_stdlogicvector(X"00");
	mem(155) := To_stdlogicvector(X"00");
	mem(156) := To_stdlogicvector(X"00");
	mem(157) := To_stdlogicvector(X"00");
	mem(158) := To_stdlogicvector(X"00");
	mem(159) := To_stdlogicvector(X"00");
	mem(160) := To_stdlogicvector(X"00");
	mem(161) := To_stdlogicvector(X"00");
	mem(162) := To_stdlogicvector(X"00");
	mem(163) := To_stdlogicvector(X"00");
	mem(164) := To_stdlogicvector(X"41");
	mem(165) := To_stdlogicvector(X"12");
	mem(166) := To_stdlogicvector(X"00");
	mem(167) := To_stdlogicvector(X"00");
	mem(168) := To_stdlogicvector(X"00");
	mem(169) := To_stdlogicvector(X"00");
	mem(170) := To_stdlogicvector(X"00");
	mem(171) := To_stdlogicvector(X"00");
	mem(172) := To_stdlogicvector(X"00");
	mem(173) := To_stdlogicvector(X"00");
	mem(174) := To_stdlogicvector(X"00");
	mem(175) := To_stdlogicvector(X"00");
	mem(176) := To_stdlogicvector(X"00");
	mem(177) := To_stdlogicvector(X"00");
	mem(178) := To_stdlogicvector(X"0F");
	mem(179) := To_stdlogicvector(X"72");
	mem(180) := To_stdlogicvector(X"00");
	mem(181) := To_stdlogicvector(X"00");
	mem(182) := To_stdlogicvector(X"00");
	mem(183) := To_stdlogicvector(X"00");
	mem(184) := To_stdlogicvector(X"00");
	mem(185) := To_stdlogicvector(X"00");
	mem(186) := To_stdlogicvector(X"00");
	mem(187) := To_stdlogicvector(X"00");
	mem(188) := To_stdlogicvector(X"00");
	mem(189) := To_stdlogicvector(X"00");
	mem(190) := To_stdlogicvector(X"00");
	mem(191) := To_stdlogicvector(X"00");
	mem(192) := To_stdlogicvector(X"03");
	mem(193) := To_stdlogicvector(X"62");
	mem(194) := To_stdlogicvector(X"00");
	mem(195) := To_stdlogicvector(X"00");
	mem(196) := To_stdlogicvector(X"00");
	mem(197) := To_stdlogicvector(X"00");
	mem(198) := To_stdlogicvector(X"00");
	mem(199) := To_stdlogicvector(X"00");
	mem(200) := To_stdlogicvector(X"00");
	mem(201) := To_stdlogicvector(X"00");
	mem(202) := To_stdlogicvector(X"00");
	mem(203) := To_stdlogicvector(X"00");
	mem(204) := To_stdlogicvector(X"00");
	mem(205) := To_stdlogicvector(X"00");
	mem(206) := To_stdlogicvector(X"04");
	mem(207) := To_stdlogicvector(X"64");
	mem(208) := To_stdlogicvector(X"00");
	mem(209) := To_stdlogicvector(X"00");
	mem(210) := To_stdlogicvector(X"00");
	mem(211) := To_stdlogicvector(X"00");
	mem(212) := To_stdlogicvector(X"00");
	mem(213) := To_stdlogicvector(X"00");
	mem(214) := To_stdlogicvector(X"00");
	mem(215) := To_stdlogicvector(X"00");
	mem(216) := To_stdlogicvector(X"00");
	mem(217) := To_stdlogicvector(X"00");
	mem(218) := To_stdlogicvector(X"00");
	mem(219) := To_stdlogicvector(X"00");
	mem(220) := To_stdlogicvector(X"42");
	mem(221) := To_stdlogicvector(X"5C");
	mem(222) := To_stdlogicvector(X"00");
	mem(223) := To_stdlogicvector(X"00");
	mem(224) := To_stdlogicvector(X"00");
	mem(225) := To_stdlogicvector(X"00");
	mem(226) := To_stdlogicvector(X"00");
	mem(227) := To_stdlogicvector(X"00");
	mem(228) := To_stdlogicvector(X"00");
	mem(229) := To_stdlogicvector(X"00");
	mem(230) := To_stdlogicvector(X"00");
	mem(231) := To_stdlogicvector(X"00");
	mem(232) := To_stdlogicvector(X"00");
	mem(233) := To_stdlogicvector(X"00");
	mem(234) := To_stdlogicvector(X"AA");
	mem(235) := To_stdlogicvector(X"5B");
	mem(236) := To_stdlogicvector(X"00");
	mem(237) := To_stdlogicvector(X"00");
	mem(238) := To_stdlogicvector(X"00");
	mem(239) := To_stdlogicvector(X"00");
	mem(240) := To_stdlogicvector(X"00");
	mem(241) := To_stdlogicvector(X"00");
	mem(242) := To_stdlogicvector(X"00");
	mem(243) := To_stdlogicvector(X"00");
	mem(244) := To_stdlogicvector(X"00");
	mem(245) := To_stdlogicvector(X"00");
	mem(246) := To_stdlogicvector(X"00");
	mem(247) := To_stdlogicvector(X"00");
	mem(248) := To_stdlogicvector(X"10");
	mem(249) := To_stdlogicvector(X"7A");
	mem(250) := To_stdlogicvector(X"00");
	mem(251) := To_stdlogicvector(X"00");
	mem(252) := To_stdlogicvector(X"00");
	mem(253) := To_stdlogicvector(X"00");
	mem(254) := To_stdlogicvector(X"00");
	mem(255) := To_stdlogicvector(X"00");
	mem(256) := To_stdlogicvector(X"00");
	mem(257) := To_stdlogicvector(X"00");
	mem(258) := To_stdlogicvector(X"00");
	mem(259) := To_stdlogicvector(X"00");
	mem(260) := To_stdlogicvector(X"00");
	mem(261) := To_stdlogicvector(X"00");
	mem(262) := To_stdlogicvector(X"05");
	mem(263) := To_stdlogicvector(X"6E");
	mem(264) := To_stdlogicvector(X"00");
	mem(265) := To_stdlogicvector(X"00");
	mem(266) := To_stdlogicvector(X"00");
	mem(267) := To_stdlogicvector(X"00");
	mem(268) := To_stdlogicvector(X"00");
	mem(269) := To_stdlogicvector(X"00");
	mem(270) := To_stdlogicvector(X"00");
	mem(271) := To_stdlogicvector(X"00");
	mem(272) := To_stdlogicvector(X"00");
	mem(273) := To_stdlogicvector(X"00");
	mem(274) := To_stdlogicvector(X"00");
	mem(275) := To_stdlogicvector(X"00");
	mem(276) := To_stdlogicvector(X"FF");
	mem(277) := To_stdlogicvector(X"9F");
	mem(278) := To_stdlogicvector(X"00");
	mem(279) := To_stdlogicvector(X"00");
	mem(280) := To_stdlogicvector(X"00");
	mem(281) := To_stdlogicvector(X"00");
	mem(282) := To_stdlogicvector(X"00");
	mem(283) := To_stdlogicvector(X"00");
	mem(284) := To_stdlogicvector(X"00");
	mem(285) := To_stdlogicvector(X"00");
	mem(286) := To_stdlogicvector(X"00");
	mem(287) := To_stdlogicvector(X"00");
	mem(288) := To_stdlogicvector(X"00");
	mem(289) := To_stdlogicvector(X"00");
	mem(290) := To_stdlogicvector(X"11");
	mem(291) := To_stdlogicvector(X"7E");
	mem(292) := To_stdlogicvector(X"00");
	mem(293) := To_stdlogicvector(X"00");
	mem(294) := To_stdlogicvector(X"00");
	mem(295) := To_stdlogicvector(X"00");
	mem(296) := To_stdlogicvector(X"00");
	mem(297) := To_stdlogicvector(X"00");
	mem(298) := To_stdlogicvector(X"00");
	mem(299) := To_stdlogicvector(X"00");
	mem(300) := To_stdlogicvector(X"00");
	mem(301) := To_stdlogicvector(X"00");
	mem(302) := To_stdlogicvector(X"00");
	mem(303) := To_stdlogicvector(X"00");
	mem(304) := To_stdlogicvector(X"09");
	mem(305) := To_stdlogicvector(X"62");
	mem(306) := To_stdlogicvector(X"00");
	mem(307) := To_stdlogicvector(X"00");
	mem(308) := To_stdlogicvector(X"00");
	mem(309) := To_stdlogicvector(X"00");
	mem(310) := To_stdlogicvector(X"00");
	mem(311) := To_stdlogicvector(X"00");
	mem(312) := To_stdlogicvector(X"00");
	mem(313) := To_stdlogicvector(X"00");
	mem(314) := To_stdlogicvector(X"00");
	mem(315) := To_stdlogicvector(X"00");
	mem(316) := To_stdlogicvector(X"00");
	mem(317) := To_stdlogicvector(X"00");
	mem(318) := To_stdlogicvector(X"64");
	mem(319) := To_stdlogicvector(X"D4");
	mem(320) := To_stdlogicvector(X"00");
	mem(321) := To_stdlogicvector(X"00");
	mem(322) := To_stdlogicvector(X"00");
	mem(323) := To_stdlogicvector(X"00");
	mem(324) := To_stdlogicvector(X"00");
	mem(325) := To_stdlogicvector(X"00");
	mem(326) := To_stdlogicvector(X"00");
	mem(327) := To_stdlogicvector(X"00");
	mem(328) := To_stdlogicvector(X"00");
	mem(329) := To_stdlogicvector(X"00");
	mem(330) := To_stdlogicvector(X"00");
	mem(331) := To_stdlogicvector(X"00");
	mem(332) := To_stdlogicvector(X"52");
	mem(333) := To_stdlogicvector(X"D6");
	mem(334) := To_stdlogicvector(X"00");
	mem(335) := To_stdlogicvector(X"00");
	mem(336) := To_stdlogicvector(X"00");
	mem(337) := To_stdlogicvector(X"00");
	mem(338) := To_stdlogicvector(X"00");
	mem(339) := To_stdlogicvector(X"00");
	mem(340) := To_stdlogicvector(X"00");
	mem(341) := To_stdlogicvector(X"00");
	mem(342) := To_stdlogicvector(X"00");
	mem(343) := To_stdlogicvector(X"00");
	mem(344) := To_stdlogicvector(X"00");
	mem(345) := To_stdlogicvector(X"00");
	mem(346) := To_stdlogicvector(X"A1");
	mem(347) := To_stdlogicvector(X"D4");
	mem(348) := To_stdlogicvector(X"00");
	mem(349) := To_stdlogicvector(X"00");
	mem(350) := To_stdlogicvector(X"00");
	mem(351) := To_stdlogicvector(X"00");
	mem(352) := To_stdlogicvector(X"00");
	mem(353) := To_stdlogicvector(X"00");
	mem(354) := To_stdlogicvector(X"00");
	mem(355) := To_stdlogicvector(X"00");
	mem(356) := To_stdlogicvector(X"00");
	mem(357) := To_stdlogicvector(X"00");
	mem(358) := To_stdlogicvector(X"00");
	mem(359) := To_stdlogicvector(X"00");
	mem(360) := To_stdlogicvector(X"D1");
	mem(361) := To_stdlogicvector(X"D6");
	mem(362) := To_stdlogicvector(X"00");
	mem(363) := To_stdlogicvector(X"00");
	mem(364) := To_stdlogicvector(X"00");
	mem(365) := To_stdlogicvector(X"00");
	mem(366) := To_stdlogicvector(X"00");
	mem(367) := To_stdlogicvector(X"00");
	mem(368) := To_stdlogicvector(X"00");
	mem(369) := To_stdlogicvector(X"00");
	mem(370) := To_stdlogicvector(X"00");
	mem(371) := To_stdlogicvector(X"00");
	mem(372) := To_stdlogicvector(X"00");
	mem(373) := To_stdlogicvector(X"00");
	mem(374) := To_stdlogicvector(X"83");
	mem(375) := To_stdlogicvector(X"14");
	mem(376) := To_stdlogicvector(X"00");
	mem(377) := To_stdlogicvector(X"00");
	mem(378) := To_stdlogicvector(X"00");
	mem(379) := To_stdlogicvector(X"00");
	mem(380) := To_stdlogicvector(X"00");
	mem(381) := To_stdlogicvector(X"00");
	mem(382) := To_stdlogicvector(X"00");
	mem(383) := To_stdlogicvector(X"00");
	mem(384) := To_stdlogicvector(X"00");
	mem(385) := To_stdlogicvector(X"00");
	mem(386) := To_stdlogicvector(X"00");
	mem(387) := To_stdlogicvector(X"00");
	mem(388) := To_stdlogicvector(X"A1");
	mem(389) := To_stdlogicvector(X"14");
	mem(390) := To_stdlogicvector(X"00");
	mem(391) := To_stdlogicvector(X"00");
	mem(392) := To_stdlogicvector(X"00");
	mem(393) := To_stdlogicvector(X"00");
	mem(394) := To_stdlogicvector(X"00");
	mem(395) := To_stdlogicvector(X"00");
	mem(396) := To_stdlogicvector(X"00");
	mem(397) := To_stdlogicvector(X"00");
	mem(398) := To_stdlogicvector(X"00");
	mem(399) := To_stdlogicvector(X"00");
	mem(400) := To_stdlogicvector(X"00");
	mem(401) := To_stdlogicvector(X"00");
	mem(402) := To_stdlogicvector(X"73");
	mem(403) := To_stdlogicvector(X"D8");
	mem(404) := To_stdlogicvector(X"00");
	mem(405) := To_stdlogicvector(X"00");
	mem(406) := To_stdlogicvector(X"00");
	mem(407) := To_stdlogicvector(X"00");
	mem(408) := To_stdlogicvector(X"00");
	mem(409) := To_stdlogicvector(X"00");
	mem(410) := To_stdlogicvector(X"00");
	mem(411) := To_stdlogicvector(X"00");
	mem(412) := To_stdlogicvector(X"00");
	mem(413) := To_stdlogicvector(X"00");
	mem(414) := To_stdlogicvector(X"00");
	mem(415) := To_stdlogicvector(X"00");
	mem(416) := To_stdlogicvector(X"0A");
	mem(417) := To_stdlogicvector(X"62");
	mem(418) := To_stdlogicvector(X"00");
	mem(419) := To_stdlogicvector(X"00");
	mem(420) := To_stdlogicvector(X"00");
	mem(421) := To_stdlogicvector(X"00");
	mem(422) := To_stdlogicvector(X"00");
	mem(423) := To_stdlogicvector(X"00");
	mem(424) := To_stdlogicvector(X"00");
	mem(425) := To_stdlogicvector(X"00");
	mem(426) := To_stdlogicvector(X"00");
	mem(427) := To_stdlogicvector(X"00");
	mem(428) := To_stdlogicvector(X"00");
	mem(429) := To_stdlogicvector(X"00");
	mem(430) := To_stdlogicvector(X"76");
	mem(431) := To_stdlogicvector(X"DA");
	mem(432) := To_stdlogicvector(X"00");
	mem(433) := To_stdlogicvector(X"00");
	mem(434) := To_stdlogicvector(X"00");
	mem(435) := To_stdlogicvector(X"00");
	mem(436) := To_stdlogicvector(X"00");
	mem(437) := To_stdlogicvector(X"00");
	mem(438) := To_stdlogicvector(X"00");
	mem(439) := To_stdlogicvector(X"00");
	mem(440) := To_stdlogicvector(X"00");
	mem(441) := To_stdlogicvector(X"00");
	mem(442) := To_stdlogicvector(X"00");
	mem(443) := To_stdlogicvector(X"00");
	mem(444) := To_stdlogicvector(X"12");
	mem(445) := To_stdlogicvector(X"74");
	mem(446) := To_stdlogicvector(X"00");
	mem(447) := To_stdlogicvector(X"00");
	mem(448) := To_stdlogicvector(X"00");
	mem(449) := To_stdlogicvector(X"00");
	mem(450) := To_stdlogicvector(X"00");
	mem(451) := To_stdlogicvector(X"00");
	mem(452) := To_stdlogicvector(X"00");
	mem(453) := To_stdlogicvector(X"00");
	mem(454) := To_stdlogicvector(X"00");
	mem(455) := To_stdlogicvector(X"00");
	mem(456) := To_stdlogicvector(X"00");
	mem(457) := To_stdlogicvector(X"00");
	mem(458) := To_stdlogicvector(X"13");
	mem(459) := To_stdlogicvector(X"78");
	mem(460) := To_stdlogicvector(X"00");
	mem(461) := To_stdlogicvector(X"00");
	mem(462) := To_stdlogicvector(X"00");
	mem(463) := To_stdlogicvector(X"00");
	mem(464) := To_stdlogicvector(X"00");
	mem(465) := To_stdlogicvector(X"00");
	mem(466) := To_stdlogicvector(X"00");
	mem(467) := To_stdlogicvector(X"00");
	mem(468) := To_stdlogicvector(X"00");
	mem(469) := To_stdlogicvector(X"00");
	mem(470) := To_stdlogicvector(X"00");
	mem(471) := To_stdlogicvector(X"00");
	mem(472) := To_stdlogicvector(X"14");
	mem(473) := To_stdlogicvector(X"7A");
	mem(474) := To_stdlogicvector(X"00");
	mem(475) := To_stdlogicvector(X"00");
	mem(476) := To_stdlogicvector(X"00");
	mem(477) := To_stdlogicvector(X"00");
	mem(478) := To_stdlogicvector(X"00");
	mem(479) := To_stdlogicvector(X"00");
	mem(480) := To_stdlogicvector(X"00");
	mem(481) := To_stdlogicvector(X"00");
	mem(482) := To_stdlogicvector(X"00");
	mem(483) := To_stdlogicvector(X"00");
	mem(484) := To_stdlogicvector(X"00");
	mem(485) := To_stdlogicvector(X"00");
	mem(486) := To_stdlogicvector(X"29");
	mem(487) := To_stdlogicvector(X"E3");
	mem(488) := To_stdlogicvector(X"00");
	mem(489) := To_stdlogicvector(X"00");
	mem(490) := To_stdlogicvector(X"00");
	mem(491) := To_stdlogicvector(X"00");
	mem(492) := To_stdlogicvector(X"00");
	mem(493) := To_stdlogicvector(X"00");
	mem(494) := To_stdlogicvector(X"00");
	mem(495) := To_stdlogicvector(X"00");
	mem(496) := To_stdlogicvector(X"00");
	mem(497) := To_stdlogicvector(X"00");
	mem(498) := To_stdlogicvector(X"00");
	mem(499) := To_stdlogicvector(X"00");
	mem(500) := To_stdlogicvector(X"16");
	mem(501) := To_stdlogicvector(X"72");
	mem(502) := To_stdlogicvector(X"00");
	mem(503) := To_stdlogicvector(X"00");
	mem(504) := To_stdlogicvector(X"00");
	mem(505) := To_stdlogicvector(X"00");
	mem(506) := To_stdlogicvector(X"00");
	mem(507) := To_stdlogicvector(X"00");
	mem(508) := To_stdlogicvector(X"00");
	mem(509) := To_stdlogicvector(X"00");
	mem(510) := To_stdlogicvector(X"00");
	mem(511) := To_stdlogicvector(X"00");
	mem(512) := To_stdlogicvector(X"00");
	mem(513) := To_stdlogicvector(X"00");
	mem(514) := To_stdlogicvector(X"6D");
	mem(515) := To_stdlogicvector(X"1B");
	mem(516) := To_stdlogicvector(X"00");
	mem(517) := To_stdlogicvector(X"00");
	mem(518) := To_stdlogicvector(X"00");
	mem(519) := To_stdlogicvector(X"00");
	mem(520) := To_stdlogicvector(X"00");
	mem(521) := To_stdlogicvector(X"00");
	mem(522) := To_stdlogicvector(X"00");
	mem(523) := To_stdlogicvector(X"00");
	mem(524) := To_stdlogicvector(X"00");
	mem(525) := To_stdlogicvector(X"00");
	mem(526) := To_stdlogicvector(X"00");
	mem(527) := To_stdlogicvector(X"00");
	mem(528) := To_stdlogicvector(X"16");
	mem(529) := To_stdlogicvector(X"BA");
	mem(530) := To_stdlogicvector(X"00");
	mem(531) := To_stdlogicvector(X"00");
	mem(532) := To_stdlogicvector(X"00");
	mem(533) := To_stdlogicvector(X"00");
	mem(534) := To_stdlogicvector(X"00");
	mem(535) := To_stdlogicvector(X"00");
	mem(536) := To_stdlogicvector(X"00");
	mem(537) := To_stdlogicvector(X"00");
	mem(538) := To_stdlogicvector(X"00");
	mem(539) := To_stdlogicvector(X"00");
	mem(540) := To_stdlogicvector(X"00");
	mem(541) := To_stdlogicvector(X"00");
	mem(542) := To_stdlogicvector(X"07");
	mem(543) := To_stdlogicvector(X"62");
	mem(544) := To_stdlogicvector(X"00");
	mem(545) := To_stdlogicvector(X"00");
	mem(546) := To_stdlogicvector(X"00");
	mem(547) := To_stdlogicvector(X"00");
	mem(548) := To_stdlogicvector(X"00");
	mem(549) := To_stdlogicvector(X"00");
	mem(550) := To_stdlogicvector(X"00");
	mem(551) := To_stdlogicvector(X"00");
	mem(552) := To_stdlogicvector(X"00");
	mem(553) := To_stdlogicvector(X"00");
	mem(554) := To_stdlogicvector(X"00");
	mem(555) := To_stdlogicvector(X"00");
	mem(556) := To_stdlogicvector(X"06");
	mem(557) := To_stdlogicvector(X"64");
	mem(558) := To_stdlogicvector(X"00");
	mem(559) := To_stdlogicvector(X"00");
	mem(560) := To_stdlogicvector(X"00");
	mem(561) := To_stdlogicvector(X"00");
	mem(562) := To_stdlogicvector(X"00");
	mem(563) := To_stdlogicvector(X"00");
	mem(564) := To_stdlogicvector(X"00");
	mem(565) := To_stdlogicvector(X"00");
	mem(566) := To_stdlogicvector(X"00");
	mem(567) := To_stdlogicvector(X"00");
	mem(568) := To_stdlogicvector(X"00");
	mem(569) := To_stdlogicvector(X"00");
	mem(570) := To_stdlogicvector(X"E0");
	mem(571) := To_stdlogicvector(X"56");
	mem(572) := To_stdlogicvector(X"00");
	mem(573) := To_stdlogicvector(X"00");
	mem(574) := To_stdlogicvector(X"00");
	mem(575) := To_stdlogicvector(X"00");
	mem(576) := To_stdlogicvector(X"00");
	mem(577) := To_stdlogicvector(X"00");
	mem(578) := To_stdlogicvector(X"00");
	mem(579) := To_stdlogicvector(X"00");
	mem(580) := To_stdlogicvector(X"00");
	mem(581) := To_stdlogicvector(X"00");
	mem(582) := To_stdlogicvector(X"00");
	mem(583) := To_stdlogicvector(X"00");
	mem(584) := To_stdlogicvector(X"A5");
	mem(585) := To_stdlogicvector(X"14");
	mem(586) := To_stdlogicvector(X"00");
	mem(587) := To_stdlogicvector(X"00");
	mem(588) := To_stdlogicvector(X"00");
	mem(589) := To_stdlogicvector(X"00");
	mem(590) := To_stdlogicvector(X"00");
	mem(591) := To_stdlogicvector(X"00");
	mem(592) := To_stdlogicvector(X"00");
	mem(593) := To_stdlogicvector(X"00");
	mem(594) := To_stdlogicvector(X"00");
	mem(595) := To_stdlogicvector(X"00");
	mem(596) := To_stdlogicvector(X"00");
	mem(597) := To_stdlogicvector(X"00");
	mem(598) := To_stdlogicvector(X"7F");
	mem(599) := To_stdlogicvector(X"12");
	mem(600) := To_stdlogicvector(X"00");
	mem(601) := To_stdlogicvector(X"00");
	mem(602) := To_stdlogicvector(X"00");
	mem(603) := To_stdlogicvector(X"00");
	mem(604) := To_stdlogicvector(X"00");
	mem(605) := To_stdlogicvector(X"00");
	mem(606) := To_stdlogicvector(X"00");
	mem(607) := To_stdlogicvector(X"00");
	mem(608) := To_stdlogicvector(X"00");
	mem(609) := To_stdlogicvector(X"00");
	mem(610) := To_stdlogicvector(X"00");
	mem(611) := To_stdlogicvector(X"00");
	mem(612) := To_stdlogicvector(X"F1");
	mem(613) := To_stdlogicvector(X"03");
	mem(614) := To_stdlogicvector(X"00");
	mem(615) := To_stdlogicvector(X"00");
	mem(616) := To_stdlogicvector(X"00");
	mem(617) := To_stdlogicvector(X"00");
	mem(618) := To_stdlogicvector(X"00");
	mem(619) := To_stdlogicvector(X"00");
	mem(620) := To_stdlogicvector(X"00");
	mem(621) := To_stdlogicvector(X"00");
	mem(622) := To_stdlogicvector(X"00");
	mem(623) := To_stdlogicvector(X"00");
	mem(624) := To_stdlogicvector(X"00");
	mem(625) := To_stdlogicvector(X"00");
	mem(626) := To_stdlogicvector(X"67");
	mem(627) := To_stdlogicvector(X"12");
	mem(628) := To_stdlogicvector(X"00");
	mem(629) := To_stdlogicvector(X"00");
	mem(630) := To_stdlogicvector(X"00");
	mem(631) := To_stdlogicvector(X"00");
	mem(632) := To_stdlogicvector(X"00");
	mem(633) := To_stdlogicvector(X"00");
	mem(634) := To_stdlogicvector(X"00");
	mem(635) := To_stdlogicvector(X"00");
	mem(636) := To_stdlogicvector(X"00");
	mem(637) := To_stdlogicvector(X"00");
	mem(638) := To_stdlogicvector(X"00");
	mem(639) := To_stdlogicvector(X"00");
	mem(640) := To_stdlogicvector(X"BA");
	mem(641) := To_stdlogicvector(X"14");
	mem(642) := To_stdlogicvector(X"00");
	mem(643) := To_stdlogicvector(X"00");
	mem(644) := To_stdlogicvector(X"00");
	mem(645) := To_stdlogicvector(X"00");
	mem(646) := To_stdlogicvector(X"00");
	mem(647) := To_stdlogicvector(X"00");
	mem(648) := To_stdlogicvector(X"00");
	mem(649) := To_stdlogicvector(X"00");
	mem(650) := To_stdlogicvector(X"00");
	mem(651) := To_stdlogicvector(X"00");
	mem(652) := To_stdlogicvector(X"00");
	mem(653) := To_stdlogicvector(X"00");
	mem(654) := To_stdlogicvector(X"F1");
	mem(655) := To_stdlogicvector(X"03");
	mem(656) := To_stdlogicvector(X"00");
	mem(657) := To_stdlogicvector(X"00");
	mem(658) := To_stdlogicvector(X"00");
	mem(659) := To_stdlogicvector(X"00");
	mem(660) := To_stdlogicvector(X"00");
	mem(661) := To_stdlogicvector(X"00");
	mem(662) := To_stdlogicvector(X"00");
	mem(663) := To_stdlogicvector(X"00");
	mem(664) := To_stdlogicvector(X"00");
	mem(665) := To_stdlogicvector(X"00");
	mem(666) := To_stdlogicvector(X"00");
	mem(667) := To_stdlogicvector(X"00");
	mem(668) := To_stdlogicvector(X"D5");
	mem(669) := To_stdlogicvector(X"05");
	mem(670) := To_stdlogicvector(X"00");
	mem(671) := To_stdlogicvector(X"00");
	mem(672) := To_stdlogicvector(X"00");
	mem(673) := To_stdlogicvector(X"00");
	mem(674) := To_stdlogicvector(X"00");
	mem(675) := To_stdlogicvector(X"00");
	mem(676) := To_stdlogicvector(X"00");
	mem(677) := To_stdlogicvector(X"00");
	mem(678) := To_stdlogicvector(X"00");
	mem(679) := To_stdlogicvector(X"00");
	mem(680) := To_stdlogicvector(X"00");
	mem(681) := To_stdlogicvector(X"00");
	mem(682) := To_stdlogicvector(X"0D");
	mem(683) := To_stdlogicvector(X"08");
	mem(684) := To_stdlogicvector(X"00");
	mem(685) := To_stdlogicvector(X"00");
	mem(686) := To_stdlogicvector(X"00");
	mem(687) := To_stdlogicvector(X"00");
	mem(688) := To_stdlogicvector(X"00");
	mem(689) := To_stdlogicvector(X"00");
	mem(690) := To_stdlogicvector(X"00");
	mem(691) := To_stdlogicvector(X"00");
	mem(692) := To_stdlogicvector(X"00");
	mem(693) := To_stdlogicvector(X"00");
	mem(694) := To_stdlogicvector(X"00");
	mem(695) := To_stdlogicvector(X"00");
	mem(696) := To_stdlogicvector(X"0D");
	mem(697) := To_stdlogicvector(X"64");
	mem(698) := To_stdlogicvector(X"00");
	mem(699) := To_stdlogicvector(X"00");
	mem(700) := To_stdlogicvector(X"00");
	mem(701) := To_stdlogicvector(X"00");
	mem(702) := To_stdlogicvector(X"00");
	mem(703) := To_stdlogicvector(X"00");
	mem(704) := To_stdlogicvector(X"00");
	mem(705) := To_stdlogicvector(X"00");
	mem(706) := To_stdlogicvector(X"00");
	mem(707) := To_stdlogicvector(X"00");
	mem(708) := To_stdlogicvector(X"00");
	mem(709) := To_stdlogicvector(X"00");
	mem(710) := To_stdlogicvector(X"81");
	mem(711) := To_stdlogicvector(X"14");
	mem(712) := To_stdlogicvector(X"00");
	mem(713) := To_stdlogicvector(X"00");
	mem(714) := To_stdlogicvector(X"00");
	mem(715) := To_stdlogicvector(X"00");
	mem(716) := To_stdlogicvector(X"00");
	mem(717) := To_stdlogicvector(X"00");
	mem(718) := To_stdlogicvector(X"00");
	mem(719) := To_stdlogicvector(X"00");
	mem(720) := To_stdlogicvector(X"00");
	mem(721) := To_stdlogicvector(X"00");
	mem(722) := To_stdlogicvector(X"00");
	mem(723) := To_stdlogicvector(X"00");
	mem(724) := To_stdlogicvector(X"16");
	mem(725) := To_stdlogicvector(X"74");
	mem(726) := To_stdlogicvector(X"00");
	mem(727) := To_stdlogicvector(X"00");
	mem(728) := To_stdlogicvector(X"00");
	mem(729) := To_stdlogicvector(X"00");
	mem(730) := To_stdlogicvector(X"00");
	mem(731) := To_stdlogicvector(X"00");
	mem(732) := To_stdlogicvector(X"00");
	mem(733) := To_stdlogicvector(X"00");
	mem(734) := To_stdlogicvector(X"00");
	mem(735) := To_stdlogicvector(X"00");
	mem(736) := To_stdlogicvector(X"00");
	mem(737) := To_stdlogicvector(X"00");
	mem(738) := To_stdlogicvector(X"00");
	mem(739) := To_stdlogicvector(X"6C");
	mem(740) := To_stdlogicvector(X"00");
	mem(741) := To_stdlogicvector(X"00");
	mem(742) := To_stdlogicvector(X"00");
	mem(743) := To_stdlogicvector(X"00");
	mem(744) := To_stdlogicvector(X"00");
	mem(745) := To_stdlogicvector(X"00");
	mem(746) := To_stdlogicvector(X"00");
	mem(747) := To_stdlogicvector(X"00");
	mem(748) := To_stdlogicvector(X"00");
	mem(749) := To_stdlogicvector(X"00");
	mem(750) := To_stdlogicvector(X"00");
	mem(751) := To_stdlogicvector(X"00");
	mem(752) := To_stdlogicvector(X"B0");
	mem(753) := To_stdlogicvector(X"49");
	mem(754) := To_stdlogicvector(X"00");
	mem(755) := To_stdlogicvector(X"00");
	mem(756) := To_stdlogicvector(X"00");
	mem(757) := To_stdlogicvector(X"00");
	mem(758) := To_stdlogicvector(X"00");
	mem(759) := To_stdlogicvector(X"00");
	mem(760) := To_stdlogicvector(X"00");
	mem(761) := To_stdlogicvector(X"00");
	mem(762) := To_stdlogicvector(X"00");
	mem(763) := To_stdlogicvector(X"00");
	mem(764) := To_stdlogicvector(X"00");
	mem(765) := To_stdlogicvector(X"00");
	mem(766) := To_stdlogicvector(X"17");
	mem(767) := To_stdlogicvector(X"7C");
	mem(768) := To_stdlogicvector(X"00");
	mem(769) := To_stdlogicvector(X"00");
	mem(770) := To_stdlogicvector(X"00");
	mem(771) := To_stdlogicvector(X"00");
	mem(772) := To_stdlogicvector(X"00");
	mem(773) := To_stdlogicvector(X"00");
	mem(774) := To_stdlogicvector(X"00");
	mem(775) := To_stdlogicvector(X"00");
	mem(776) := To_stdlogicvector(X"00");
	mem(777) := To_stdlogicvector(X"00");
	mem(778) := To_stdlogicvector(X"00");
	mem(779) := To_stdlogicvector(X"00");
	mem(780) := To_stdlogicvector(X"6D");
	mem(781) := To_stdlogicvector(X"5B");
	mem(782) := To_stdlogicvector(X"00");
	mem(783) := To_stdlogicvector(X"00");
	mem(784) := To_stdlogicvector(X"00");
	mem(785) := To_stdlogicvector(X"00");
	mem(786) := To_stdlogicvector(X"00");
	mem(787) := To_stdlogicvector(X"00");
	mem(788) := To_stdlogicvector(X"00");
	mem(789) := To_stdlogicvector(X"00");
	mem(790) := To_stdlogicvector(X"00");
	mem(791) := To_stdlogicvector(X"00");
	mem(792) := To_stdlogicvector(X"00");
	mem(793) := To_stdlogicvector(X"00");
	mem(794) := To_stdlogicvector(X"14");
	mem(795) := To_stdlogicvector(X"E6");
	mem(796) := To_stdlogicvector(X"00");
	mem(797) := To_stdlogicvector(X"00");
	mem(798) := To_stdlogicvector(X"00");
	mem(799) := To_stdlogicvector(X"00");
	mem(800) := To_stdlogicvector(X"00");
	mem(801) := To_stdlogicvector(X"00");
	mem(802) := To_stdlogicvector(X"00");
	mem(803) := To_stdlogicvector(X"00");
	mem(804) := To_stdlogicvector(X"00");
	mem(805) := To_stdlogicvector(X"00");
	mem(806) := To_stdlogicvector(X"00");
	mem(807) := To_stdlogicvector(X"00");
	mem(808) := To_stdlogicvector(X"C0");
	mem(809) := To_stdlogicvector(X"C0");
	mem(810) := To_stdlogicvector(X"00");
	mem(811) := To_stdlogicvector(X"00");
	mem(812) := To_stdlogicvector(X"00");
	mem(813) := To_stdlogicvector(X"00");
	mem(814) := To_stdlogicvector(X"00");
	mem(815) := To_stdlogicvector(X"00");
	mem(816) := To_stdlogicvector(X"00");
	mem(817) := To_stdlogicvector(X"00");
	mem(818) := To_stdlogicvector(X"00");
	mem(819) := To_stdlogicvector(X"00");
	mem(820) := To_stdlogicvector(X"00");
	mem(821) := To_stdlogicvector(X"00");
	mem(822) := To_stdlogicvector(X"08");
	mem(823) := To_stdlogicvector(X"6A");
	mem(824) := To_stdlogicvector(X"00");
	mem(825) := To_stdlogicvector(X"00");
	mem(826) := To_stdlogicvector(X"00");
	mem(827) := To_stdlogicvector(X"00");
	mem(828) := To_stdlogicvector(X"00");
	mem(829) := To_stdlogicvector(X"00");
	mem(830) := To_stdlogicvector(X"00");
	mem(831) := To_stdlogicvector(X"00");
	mem(832) := To_stdlogicvector(X"00");
	mem(833) := To_stdlogicvector(X"00");
	mem(834) := To_stdlogicvector(X"00");
	mem(835) := To_stdlogicvector(X"00");
	mem(836) := To_stdlogicvector(X"18");
	mem(837) := To_stdlogicvector(X"7A");
	mem(838) := To_stdlogicvector(X"00");
	mem(839) := To_stdlogicvector(X"00");
	mem(840) := To_stdlogicvector(X"00");
	mem(841) := To_stdlogicvector(X"00");
	mem(842) := To_stdlogicvector(X"00");
	mem(843) := To_stdlogicvector(X"00");
	mem(844) := To_stdlogicvector(X"00");
	mem(845) := To_stdlogicvector(X"00");
	mem(846) := To_stdlogicvector(X"00");
	mem(847) := To_stdlogicvector(X"00");
	mem(848) := To_stdlogicvector(X"00");
	mem(849) := To_stdlogicvector(X"00");
	mem(850) := To_stdlogicvector(X"08");
	mem(851) := To_stdlogicvector(X"6A");
	mem(852) := To_stdlogicvector(X"00");
	mem(853) := To_stdlogicvector(X"00");
	mem(854) := To_stdlogicvector(X"00");
	mem(855) := To_stdlogicvector(X"00");
	mem(856) := To_stdlogicvector(X"00");
	mem(857) := To_stdlogicvector(X"00");
	mem(858) := To_stdlogicvector(X"00");
	mem(859) := To_stdlogicvector(X"00");
	mem(860) := To_stdlogicvector(X"00");
	mem(861) := To_stdlogicvector(X"00");
	mem(862) := To_stdlogicvector(X"00");
	mem(863) := To_stdlogicvector(X"00");
	mem(864) := To_stdlogicvector(X"27");
	mem(865) := To_stdlogicvector(X"F0");
	mem(866) := To_stdlogicvector(X"00");
	mem(867) := To_stdlogicvector(X"00");
	mem(868) := To_stdlogicvector(X"00");
	mem(869) := To_stdlogicvector(X"00");
	mem(870) := To_stdlogicvector(X"00");
	mem(871) := To_stdlogicvector(X"00");
	mem(872) := To_stdlogicvector(X"00");
	mem(873) := To_stdlogicvector(X"00");
	mem(874) := To_stdlogicvector(X"00");
	mem(875) := To_stdlogicvector(X"00");
	mem(876) := To_stdlogicvector(X"00");
	mem(877) := To_stdlogicvector(X"00");
	mem(878) := To_stdlogicvector(X"19");
	mem(879) := To_stdlogicvector(X"7A");
	mem(880) := To_stdlogicvector(X"00");
	mem(881) := To_stdlogicvector(X"00");
	mem(882) := To_stdlogicvector(X"00");
	mem(883) := To_stdlogicvector(X"00");
	mem(884) := To_stdlogicvector(X"00");
	mem(885) := To_stdlogicvector(X"00");
	mem(886) := To_stdlogicvector(X"00");
	mem(887) := To_stdlogicvector(X"00");
	mem(888) := To_stdlogicvector(X"00");
	mem(889) := To_stdlogicvector(X"00");
	mem(890) := To_stdlogicvector(X"00");
	mem(891) := To_stdlogicvector(X"00");
	mem(892) := To_stdlogicvector(X"60");
	mem(893) := To_stdlogicvector(X"52");
	mem(894) := To_stdlogicvector(X"00");
	mem(895) := To_stdlogicvector(X"00");
	mem(896) := To_stdlogicvector(X"00");
	mem(897) := To_stdlogicvector(X"00");
	mem(898) := To_stdlogicvector(X"00");
	mem(899) := To_stdlogicvector(X"00");
	mem(900) := To_stdlogicvector(X"00");
	mem(901) := To_stdlogicvector(X"00");
	mem(902) := To_stdlogicvector(X"00");
	mem(903) := To_stdlogicvector(X"00");
	mem(904) := To_stdlogicvector(X"00");
	mem(905) := To_stdlogicvector(X"00");
	mem(906) := To_stdlogicvector(X"68");
	mem(907) := To_stdlogicvector(X"12");
	mem(908) := To_stdlogicvector(X"00");
	mem(909) := To_stdlogicvector(X"00");
	mem(910) := To_stdlogicvector(X"00");
	mem(911) := To_stdlogicvector(X"00");
	mem(912) := To_stdlogicvector(X"00");
	mem(913) := To_stdlogicvector(X"00");
	mem(914) := To_stdlogicvector(X"00");
	mem(915) := To_stdlogicvector(X"00");
	mem(916) := To_stdlogicvector(X"00");
	mem(917) := To_stdlogicvector(X"00");
	mem(918) := To_stdlogicvector(X"00");
	mem(919) := To_stdlogicvector(X"00");
	mem(920) := To_stdlogicvector(X"69");
	mem(921) := To_stdlogicvector(X"12");
	mem(922) := To_stdlogicvector(X"00");
	mem(923) := To_stdlogicvector(X"00");
	mem(924) := To_stdlogicvector(X"00");
	mem(925) := To_stdlogicvector(X"00");
	mem(926) := To_stdlogicvector(X"00");
	mem(927) := To_stdlogicvector(X"00");
	mem(928) := To_stdlogicvector(X"00");
	mem(929) := To_stdlogicvector(X"00");
	mem(930) := To_stdlogicvector(X"00");
	mem(931) := To_stdlogicvector(X"00");
	mem(932) := To_stdlogicvector(X"00");
	mem(933) := To_stdlogicvector(X"00");
	mem(934) := To_stdlogicvector(X"16");
	mem(935) := To_stdlogicvector(X"24");
	mem(936) := To_stdlogicvector(X"00");
	mem(937) := To_stdlogicvector(X"00");
	mem(938) := To_stdlogicvector(X"00");
	mem(939) := To_stdlogicvector(X"00");
	mem(940) := To_stdlogicvector(X"00");
	mem(941) := To_stdlogicvector(X"00");
	mem(942) := To_stdlogicvector(X"00");
	mem(943) := To_stdlogicvector(X"00");
	mem(944) := To_stdlogicvector(X"00");
	mem(945) := To_stdlogicvector(X"00");
	mem(946) := To_stdlogicvector(X"00");
	mem(947) := To_stdlogicvector(X"00");
	mem(948) := To_stdlogicvector(X"56");
	mem(949) := To_stdlogicvector(X"26");
	mem(950) := To_stdlogicvector(X"00");
	mem(951) := To_stdlogicvector(X"00");
	mem(952) := To_stdlogicvector(X"00");
	mem(953) := To_stdlogicvector(X"00");
	mem(954) := To_stdlogicvector(X"00");
	mem(955) := To_stdlogicvector(X"00");
	mem(956) := To_stdlogicvector(X"00");
	mem(957) := To_stdlogicvector(X"00");
	mem(958) := To_stdlogicvector(X"00");
	mem(959) := To_stdlogicvector(X"00");
	mem(960) := To_stdlogicvector(X"00");
	mem(961) := To_stdlogicvector(X"00");
	mem(962) := To_stdlogicvector(X"C2");
	mem(963) := To_stdlogicvector(X"18");
	mem(964) := To_stdlogicvector(X"00");
	mem(965) := To_stdlogicvector(X"00");
	mem(966) := To_stdlogicvector(X"00");
	mem(967) := To_stdlogicvector(X"00");
	mem(968) := To_stdlogicvector(X"00");
	mem(969) := To_stdlogicvector(X"00");
	mem(970) := To_stdlogicvector(X"00");
	mem(971) := To_stdlogicvector(X"00");
	mem(972) := To_stdlogicvector(X"00");
	mem(973) := To_stdlogicvector(X"00");
	mem(974) := To_stdlogicvector(X"00");
	mem(975) := To_stdlogicvector(X"00");
	mem(976) := To_stdlogicvector(X"1A");
	mem(977) := To_stdlogicvector(X"78");
	mem(978) := To_stdlogicvector(X"00");
	mem(979) := To_stdlogicvector(X"00");
	mem(980) := To_stdlogicvector(X"00");
	mem(981) := To_stdlogicvector(X"00");
	mem(982) := To_stdlogicvector(X"00");
	mem(983) := To_stdlogicvector(X"00");
	mem(984) := To_stdlogicvector(X"00");
	mem(985) := To_stdlogicvector(X"00");
	mem(986) := To_stdlogicvector(X"00");
	mem(987) := To_stdlogicvector(X"00");
	mem(988) := To_stdlogicvector(X"00");
	mem(989) := To_stdlogicvector(X"00");
	mem(990) := To_stdlogicvector(X"AB");
	mem(991) := To_stdlogicvector(X"14");
	mem(992) := To_stdlogicvector(X"00");
	mem(993) := To_stdlogicvector(X"00");
	mem(994) := To_stdlogicvector(X"00");
	mem(995) := To_stdlogicvector(X"00");
	mem(996) := To_stdlogicvector(X"00");
	mem(997) := To_stdlogicvector(X"00");
	mem(998) := To_stdlogicvector(X"00");
	mem(999) := To_stdlogicvector(X"00");
	mem(1000) := To_stdlogicvector(X"00");
	mem(1001) := To_stdlogicvector(X"00");
	mem(1002) := To_stdlogicvector(X"00");
	mem(1003) := To_stdlogicvector(X"00");
	mem(1004) := To_stdlogicvector(X"FE");
	mem(1005) := To_stdlogicvector(X"16");
	mem(1006) := To_stdlogicvector(X"00");
	mem(1007) := To_stdlogicvector(X"00");
	mem(1008) := To_stdlogicvector(X"00");
	mem(1009) := To_stdlogicvector(X"00");
	mem(1010) := To_stdlogicvector(X"00");
	mem(1011) := To_stdlogicvector(X"00");
	mem(1012) := To_stdlogicvector(X"00");
	mem(1013) := To_stdlogicvector(X"00");
	mem(1014) := To_stdlogicvector(X"00");
	mem(1015) := To_stdlogicvector(X"00");
	mem(1016) := To_stdlogicvector(X"00");
	mem(1017) := To_stdlogicvector(X"00");
	mem(1018) := To_stdlogicvector(X"0D");
	mem(1019) := To_stdlogicvector(X"E2");
	mem(1020) := To_stdlogicvector(X"00");
	mem(1021) := To_stdlogicvector(X"00");
	mem(1022) := To_stdlogicvector(X"00");
	mem(1023) := To_stdlogicvector(X"00");
	mem(1024) := To_stdlogicvector(X"00");
	mem(1025) := To_stdlogicvector(X"00");
	mem(1026) := To_stdlogicvector(X"00");
	mem(1027) := To_stdlogicvector(X"00");
	mem(1028) := To_stdlogicvector(X"00");
	mem(1029) := To_stdlogicvector(X"00");
	mem(1030) := To_stdlogicvector(X"00");
	mem(1031) := To_stdlogicvector(X"00");
	mem(1032) := To_stdlogicvector(X"34");
	mem(1033) := To_stdlogicvector(X"0E");
	mem(1034) := To_stdlogicvector(X"00");
	mem(1035) := To_stdlogicvector(X"00");
	mem(1036) := To_stdlogicvector(X"00");
	mem(1037) := To_stdlogicvector(X"00");
	mem(1038) := To_stdlogicvector(X"00");
	mem(1039) := To_stdlogicvector(X"00");
	mem(1040) := To_stdlogicvector(X"00");
	mem(1041) := To_stdlogicvector(X"00");
	mem(1042) := To_stdlogicvector(X"00");
	mem(1043) := To_stdlogicvector(X"00");
	mem(1044) := To_stdlogicvector(X"00");
	mem(1045) := To_stdlogicvector(X"00");
	mem(1046) := To_stdlogicvector(X"46");
	mem(1047) := To_stdlogicvector(X"06");
	mem(1048) := To_stdlogicvector(X"00");
	mem(1049) := To_stdlogicvector(X"00");
	mem(1050) := To_stdlogicvector(X"00");
	mem(1051) := To_stdlogicvector(X"00");
	mem(1052) := To_stdlogicvector(X"00");
	mem(1053) := To_stdlogicvector(X"00");
	mem(1054) := To_stdlogicvector(X"0B");
	mem(1055) := To_stdlogicvector(X"6A");
	mem(1056) := To_stdlogicvector(X"00");
	mem(1057) := To_stdlogicvector(X"00");
	mem(1058) := To_stdlogicvector(X"00");
	mem(1059) := To_stdlogicvector(X"00");
	mem(1060) := To_stdlogicvector(X"00");
	mem(1061) := To_stdlogicvector(X"00");
	mem(1062) := To_stdlogicvector(X"00");
	mem(1063) := To_stdlogicvector(X"00");
	mem(1064) := To_stdlogicvector(X"00");
	mem(1065) := To_stdlogicvector(X"00");
	mem(1066) := To_stdlogicvector(X"00");
	mem(1067) := To_stdlogicvector(X"00");
	mem(1068) := To_stdlogicvector(X"7F");
	mem(1069) := To_stdlogicvector(X"9B");
	mem(1070) := To_stdlogicvector(X"00");
	mem(1071) := To_stdlogicvector(X"00");
	mem(1072) := To_stdlogicvector(X"00");
	mem(1073) := To_stdlogicvector(X"00");
	mem(1074) := To_stdlogicvector(X"00");
	mem(1075) := To_stdlogicvector(X"00");
	mem(1076) := To_stdlogicvector(X"00");
	mem(1077) := To_stdlogicvector(X"00");
	mem(1078) := To_stdlogicvector(X"00");
	mem(1079) := To_stdlogicvector(X"00");
	mem(1080) := To_stdlogicvector(X"00");
	mem(1081) := To_stdlogicvector(X"00");
	mem(1082) := To_stdlogicvector(X"C0");
	mem(1083) := To_stdlogicvector(X"C1");
	mem(1084) := To_stdlogicvector(X"00");
	mem(1085) := To_stdlogicvector(X"00");
	mem(1086) := To_stdlogicvector(X"00");
	mem(1087) := To_stdlogicvector(X"00");
	mem(1088) := To_stdlogicvector(X"00");
	mem(1089) := To_stdlogicvector(X"00");
	mem(1090) := To_stdlogicvector(X"00");
	mem(1091) := To_stdlogicvector(X"00");
	mem(1092) := To_stdlogicvector(X"00");
	mem(1093) := To_stdlogicvector(X"00");
	mem(1094) := To_stdlogicvector(X"00");
	mem(1095) := To_stdlogicvector(X"00");
	mem(1096) := To_stdlogicvector(X"0C");
	mem(1097) := To_stdlogicvector(X"66");
	mem(1098) := To_stdlogicvector(X"00");
	mem(1099) := To_stdlogicvector(X"00");
	mem(1100) := To_stdlogicvector(X"00");
	mem(1101) := To_stdlogicvector(X"00");
	mem(1102) := To_stdlogicvector(X"00");
	mem(1103) := To_stdlogicvector(X"00");
	mem(1104) := To_stdlogicvector(X"00");
	mem(1105) := To_stdlogicvector(X"00");
	mem(1106) := To_stdlogicvector(X"00");
	mem(1107) := To_stdlogicvector(X"00");
	mem(1108) := To_stdlogicvector(X"00");
	mem(1109) := To_stdlogicvector(X"00");
	mem(1110) := To_stdlogicvector(X"43");
	mem(1111) := To_stdlogicvector(X"12");
	mem(1112) := To_stdlogicvector(X"00");
	mem(1113) := To_stdlogicvector(X"00");
	mem(1114) := To_stdlogicvector(X"00");
	mem(1115) := To_stdlogicvector(X"00");
	mem(1116) := To_stdlogicvector(X"00");
	mem(1117) := To_stdlogicvector(X"00");
	mem(1118) := To_stdlogicvector(X"00");
	mem(1119) := To_stdlogicvector(X"00");
	mem(1120) := To_stdlogicvector(X"00");
	mem(1121) := To_stdlogicvector(X"00");
	mem(1122) := To_stdlogicvector(X"00");
	mem(1123) := To_stdlogicvector(X"00");
	mem(1124) := To_stdlogicvector(X"C0");
	mem(1125) := To_stdlogicvector(X"C1");
	mem(1126) := To_stdlogicvector(X"00");
	mem(1127) := To_stdlogicvector(X"00");
	mem(1128) := To_stdlogicvector(X"00");
	mem(1129) := To_stdlogicvector(X"00");
	mem(1130) := To_stdlogicvector(X"00");
	mem(1131) := To_stdlogicvector(X"00");
	mem(1132) := To_stdlogicvector(X"00");
	mem(1133) := To_stdlogicvector(X"00");
	mem(1134) := To_stdlogicvector(X"00");
	mem(1135) := To_stdlogicvector(X"00");
	mem(1136) := To_stdlogicvector(X"00");
	mem(1137) := To_stdlogicvector(X"00");
	mem(1138) := To_stdlogicvector(X"43");
	mem(1139) := To_stdlogicvector(X"34");
	mem(1140) := To_stdlogicvector(X"00");
	mem(1141) := To_stdlogicvector(X"00");
	mem(1142) := To_stdlogicvector(X"00");
	mem(1143) := To_stdlogicvector(X"00");
	mem(1144) := To_stdlogicvector(X"00");
	mem(1145) := To_stdlogicvector(X"00");
	mem(1146) := To_stdlogicvector(X"00");
	mem(1147) := To_stdlogicvector(X"00");
	mem(1148) := To_stdlogicvector(X"00");
	mem(1149) := To_stdlogicvector(X"00");
	mem(1150) := To_stdlogicvector(X"00");
	mem(1151) := To_stdlogicvector(X"00");
	mem(1152) := To_stdlogicvector(X"42");
	mem(1153) := To_stdlogicvector(X"36");
	mem(1154) := To_stdlogicvector(X"00");
	mem(1155) := To_stdlogicvector(X"00");
	mem(1156) := To_stdlogicvector(X"00");
	mem(1157) := To_stdlogicvector(X"00");
	mem(1158) := To_stdlogicvector(X"00");
	mem(1159) := To_stdlogicvector(X"00");
	mem(1160) := To_stdlogicvector(X"00");
	mem(1161) := To_stdlogicvector(X"00");
	mem(1162) := To_stdlogicvector(X"00");
	mem(1163) := To_stdlogicvector(X"00");
	mem(1164) := To_stdlogicvector(X"00");
	mem(1165) := To_stdlogicvector(X"00");
	mem(1166) := To_stdlogicvector(X"41");
	mem(1167) := To_stdlogicvector(X"68");
	mem(1168) := To_stdlogicvector(X"00");
	mem(1169) := To_stdlogicvector(X"00");
	mem(1170) := To_stdlogicvector(X"00");
	mem(1171) := To_stdlogicvector(X"00");
	mem(1172) := To_stdlogicvector(X"00");
	mem(1173) := To_stdlogicvector(X"00");
	mem(1174) := To_stdlogicvector(X"00");
	mem(1175) := To_stdlogicvector(X"00");
	mem(1176) := To_stdlogicvector(X"00");
	mem(1177) := To_stdlogicvector(X"00");
	mem(1178) := To_stdlogicvector(X"00");
	mem(1179) := To_stdlogicvector(X"00");
	mem(1180) := To_stdlogicvector(X"1A");
	mem(1181) := To_stdlogicvector(X"78");
	mem(1182) := To_stdlogicvector(X"00");
	mem(1183) := To_stdlogicvector(X"00");
	mem(1184) := To_stdlogicvector(X"00");
	mem(1185) := To_stdlogicvector(X"00");
	mem(1186) := To_stdlogicvector(X"00");
	mem(1187) := To_stdlogicvector(X"00");
	mem(1188) := To_stdlogicvector(X"00");
	mem(1189) := To_stdlogicvector(X"00");
	mem(1190) := To_stdlogicvector(X"00");
	mem(1191) := To_stdlogicvector(X"00");
	mem(1192) := To_stdlogicvector(X"00");
	mem(1193) := To_stdlogicvector(X"00");
	mem(1194) := To_stdlogicvector(X"B5");
	mem(1195) := To_stdlogicvector(X"E7");
	mem(1196) := To_stdlogicvector(X"00");
	mem(1197) := To_stdlogicvector(X"00");
	mem(1198) := To_stdlogicvector(X"00");
	mem(1199) := To_stdlogicvector(X"00");
	mem(1200) := To_stdlogicvector(X"00");
	mem(1201) := To_stdlogicvector(X"00");
	mem(1202) := To_stdlogicvector(X"00");
	mem(1203) := To_stdlogicvector(X"00");
	mem(1204) := To_stdlogicvector(X"00");
	mem(1205) := To_stdlogicvector(X"00");
	mem(1206) := To_stdlogicvector(X"00");
	mem(1207) := To_stdlogicvector(X"00");
	mem(1208) := To_stdlogicvector(X"1D");
	mem(1209) := To_stdlogicvector(X"76");
	mem(1210) := To_stdlogicvector(X"00");
	mem(1211) := To_stdlogicvector(X"00");
	mem(1212) := To_stdlogicvector(X"00");
	mem(1213) := To_stdlogicvector(X"00");
	mem(1214) := To_stdlogicvector(X"00");
	mem(1215) := To_stdlogicvector(X"00");
	mem(1216) := To_stdlogicvector(X"00");
	mem(1217) := To_stdlogicvector(X"00");
	mem(1218) := To_stdlogicvector(X"00");
	mem(1219) := To_stdlogicvector(X"00");
	mem(1220) := To_stdlogicvector(X"00");
	mem(1221) := To_stdlogicvector(X"00");
	mem(1222) := To_stdlogicvector(X"1D");
	mem(1223) := To_stdlogicvector(X"A6");
	mem(1224) := To_stdlogicvector(X"00");
	mem(1225) := To_stdlogicvector(X"00");
	mem(1226) := To_stdlogicvector(X"00");
	mem(1227) := To_stdlogicvector(X"00");
	mem(1228) := To_stdlogicvector(X"00");
	mem(1229) := To_stdlogicvector(X"00");
	mem(1230) := To_stdlogicvector(X"00");
	mem(1231) := To_stdlogicvector(X"00");
	mem(1232) := To_stdlogicvector(X"00");
	mem(1233) := To_stdlogicvector(X"00");
	mem(1234) := To_stdlogicvector(X"00");
	mem(1235) := To_stdlogicvector(X"00");
	mem(1236) := To_stdlogicvector(X"1C");
	mem(1237) := To_stdlogicvector(X"76");
	mem(1238) := To_stdlogicvector(X"00");
	mem(1239) := To_stdlogicvector(X"00");
	mem(1240) := To_stdlogicvector(X"00");
	mem(1241) := To_stdlogicvector(X"00");
	mem(1242) := To_stdlogicvector(X"00");
	mem(1243) := To_stdlogicvector(X"00");
	mem(1244) := To_stdlogicvector(X"00");
	mem(1245) := To_stdlogicvector(X"00");
	mem(1246) := To_stdlogicvector(X"00");
	mem(1247) := To_stdlogicvector(X"00");
	mem(1248) := To_stdlogicvector(X"00");
	mem(1249) := To_stdlogicvector(X"00");
	mem(1250) := To_stdlogicvector(X"1B");
	mem(1251) := To_stdlogicvector(X"E8");
	mem(1252) := To_stdlogicvector(X"00");
	mem(1253) := To_stdlogicvector(X"00");
	mem(1254) := To_stdlogicvector(X"00");
	mem(1255) := To_stdlogicvector(X"00");
	mem(1256) := To_stdlogicvector(X"00");
	mem(1257) := To_stdlogicvector(X"00");
	mem(1258) := To_stdlogicvector(X"00");
	mem(1259) := To_stdlogicvector(X"00");
	mem(1260) := To_stdlogicvector(X"00");
	mem(1261) := To_stdlogicvector(X"00");
	mem(1262) := To_stdlogicvector(X"00");
	mem(1263) := To_stdlogicvector(X"00");
	mem(1264) := To_stdlogicvector(X"00");
	mem(1265) := To_stdlogicvector(X"65");
	mem(1266) := To_stdlogicvector(X"00");
	mem(1267) := To_stdlogicvector(X"00");
	mem(1268) := To_stdlogicvector(X"00");
	mem(1269) := To_stdlogicvector(X"00");
	mem(1270) := To_stdlogicvector(X"00");
	mem(1271) := To_stdlogicvector(X"00");
	mem(1272) := To_stdlogicvector(X"00");
	mem(1273) := To_stdlogicvector(X"00");
	mem(1274) := To_stdlogicvector(X"00");
	mem(1275) := To_stdlogicvector(X"00");
	mem(1276) := To_stdlogicvector(X"00");
	mem(1277) := To_stdlogicvector(X"00");
	mem(1278) := To_stdlogicvector(X"A3");
	mem(1279) := To_stdlogicvector(X"14");
	mem(1280) := To_stdlogicvector(X"00");
	mem(1281) := To_stdlogicvector(X"00");
	mem(1282) := To_stdlogicvector(X"00");
	mem(1283) := To_stdlogicvector(X"00");
	mem(1284) := To_stdlogicvector(X"00");
	mem(1285) := To_stdlogicvector(X"00");
	mem(1286) := To_stdlogicvector(X"00");
	mem(1287) := To_stdlogicvector(X"00");
	mem(1288) := To_stdlogicvector(X"00");
	mem(1289) := To_stdlogicvector(X"00");
	mem(1290) := To_stdlogicvector(X"00");
	mem(1291) := To_stdlogicvector(X"00");
	mem(1292) := To_stdlogicvector(X"60");
	mem(1293) := To_stdlogicvector(X"52");
	mem(1294) := To_stdlogicvector(X"00");
	mem(1295) := To_stdlogicvector(X"00");
	mem(1296) := To_stdlogicvector(X"00");
	mem(1297) := To_stdlogicvector(X"00");
	mem(1298) := To_stdlogicvector(X"00");
	mem(1299) := To_stdlogicvector(X"00");
	mem(1300) := To_stdlogicvector(X"00");
	mem(1301) := To_stdlogicvector(X"00");
	mem(1302) := To_stdlogicvector(X"00");
	mem(1303) := To_stdlogicvector(X"00");
	mem(1304) := To_stdlogicvector(X"00");
	mem(1305) := To_stdlogicvector(X"00");
	mem(1306) := To_stdlogicvector(X"6C");
	mem(1307) := To_stdlogicvector(X"12");
	mem(1308) := To_stdlogicvector(X"00");
	mem(1309) := To_stdlogicvector(X"00");
	mem(1310) := To_stdlogicvector(X"00");
	mem(1311) := To_stdlogicvector(X"00");
	mem(1312) := To_stdlogicvector(X"00");
	mem(1313) := To_stdlogicvector(X"00");
	mem(1314) := To_stdlogicvector(X"00");
	mem(1315) := To_stdlogicvector(X"00");
	mem(1316) := To_stdlogicvector(X"00");
	mem(1317) := To_stdlogicvector(X"00");
	mem(1318) := To_stdlogicvector(X"00");
	mem(1319) := To_stdlogicvector(X"00");
	mem(1320) := To_stdlogicvector(X"1E");
	mem(1321) := To_stdlogicvector(X"72");
	mem(1322) := To_stdlogicvector(X"00");
	mem(1323) := To_stdlogicvector(X"00");
	mem(1324) := To_stdlogicvector(X"00");
	mem(1325) := To_stdlogicvector(X"00");
	mem(1326) := To_stdlogicvector(X"00");
	mem(1327) := To_stdlogicvector(X"00");
	mem(1328) := To_stdlogicvector(X"00");
	mem(1329) := To_stdlogicvector(X"00");
	mem(1330) := To_stdlogicvector(X"00");
	mem(1331) := To_stdlogicvector(X"00");
	mem(1332) := To_stdlogicvector(X"00");
	mem(1333) := To_stdlogicvector(X"00");
	mem(1334) := To_stdlogicvector(X"21");
	mem(1335) := To_stdlogicvector(X"12");
	mem(1336) := To_stdlogicvector(X"00");
	mem(1337) := To_stdlogicvector(X"00");
	mem(1338) := To_stdlogicvector(X"00");
	mem(1339) := To_stdlogicvector(X"00");
	mem(1340) := To_stdlogicvector(X"00");
	mem(1341) := To_stdlogicvector(X"00");
	mem(1342) := To_stdlogicvector(X"00");
	mem(1343) := To_stdlogicvector(X"00");
	mem(1344) := To_stdlogicvector(X"00");
	mem(1345) := To_stdlogicvector(X"00");
	mem(1346) := To_stdlogicvector(X"00");
	mem(1347) := To_stdlogicvector(X"00");
	mem(1348) := To_stdlogicvector(X"4B");
	mem(1349) := To_stdlogicvector(X"66");
	mem(1350) := To_stdlogicvector(X"00");
	mem(1351) := To_stdlogicvector(X"00");
	mem(1352) := To_stdlogicvector(X"00");
	mem(1353) := To_stdlogicvector(X"00");
	mem(1354) := To_stdlogicvector(X"00");
	mem(1355) := To_stdlogicvector(X"00");
	mem(1356) := To_stdlogicvector(X"00");
	mem(1357) := To_stdlogicvector(X"00");
	mem(1358) := To_stdlogicvector(X"00");
	mem(1359) := To_stdlogicvector(X"00");
	mem(1360) := To_stdlogicvector(X"00");
	mem(1361) := To_stdlogicvector(X"00");
	mem(1362) := To_stdlogicvector(X"61");
	mem(1363) := To_stdlogicvector(X"ED");
	mem(1364) := To_stdlogicvector(X"00");
	mem(1365) := To_stdlogicvector(X"00");
	mem(1366) := To_stdlogicvector(X"00");
	mem(1367) := To_stdlogicvector(X"00");
	mem(1368) := To_stdlogicvector(X"00");
	mem(1369) := To_stdlogicvector(X"00");
	mem(1370) := To_stdlogicvector(X"00");
	mem(1371) := To_stdlogicvector(X"00");
	mem(1372) := To_stdlogicvector(X"00");
	mem(1373) := To_stdlogicvector(X"00");
	mem(1374) := To_stdlogicvector(X"00");
	mem(1375) := To_stdlogicvector(X"00");
	mem(1376) := To_stdlogicvector(X"81");
	mem(1377) := To_stdlogicvector(X"77");
	mem(1378) := To_stdlogicvector(X"00");
	mem(1379) := To_stdlogicvector(X"00");
	mem(1380) := To_stdlogicvector(X"00");
	mem(1381) := To_stdlogicvector(X"00");
	mem(1382) := To_stdlogicvector(X"00");
	mem(1383) := To_stdlogicvector(X"00");
	mem(1384) := To_stdlogicvector(X"00");
	mem(1385) := To_stdlogicvector(X"00");
	mem(1386) := To_stdlogicvector(X"00");
	mem(1387) := To_stdlogicvector(X"00");
	mem(1388) := To_stdlogicvector(X"00");
	mem(1389) := To_stdlogicvector(X"00");
	mem(1390) := To_stdlogicvector(X"0B");
	mem(1391) := To_stdlogicvector(X"62");
	mem(1392) := To_stdlogicvector(X"00");
	mem(1393) := To_stdlogicvector(X"00");
	mem(1394) := To_stdlogicvector(X"00");
	mem(1395) := To_stdlogicvector(X"00");
	mem(1396) := To_stdlogicvector(X"00");
	mem(1397) := To_stdlogicvector(X"00");
	mem(1398) := To_stdlogicvector(X"00");
	mem(1399) := To_stdlogicvector(X"00");
	mem(1400) := To_stdlogicvector(X"00");
	mem(1401) := To_stdlogicvector(X"00");
	mem(1402) := To_stdlogicvector(X"00");
	mem(1403) := To_stdlogicvector(X"00");
	mem(1404) := To_stdlogicvector(X"78");
	mem(1405) := To_stdlogicvector(X"06");
	mem(1406) := To_stdlogicvector(X"00");
	mem(1407) := To_stdlogicvector(X"00");
	mem(1408) := To_stdlogicvector(X"00");
	mem(1409) := To_stdlogicvector(X"00");
	mem(1410) := To_stdlogicvector(X"00");
	mem(1411) := To_stdlogicvector(X"00");
	mem(1412) := To_stdlogicvector(X"00");
	mem(1413) := To_stdlogicvector(X"00");
	mem(1414) := To_stdlogicvector(X"00");
	mem(1415) := To_stdlogicvector(X"00");
	mem(1416) := To_stdlogicvector(X"00");
	mem(1417) := To_stdlogicvector(X"00");
	mem(1418) := To_stdlogicvector(X"08");
	mem(1419) := To_stdlogicvector(X"62");
	mem(1420) := To_stdlogicvector(X"00");
	mem(1421) := To_stdlogicvector(X"00");
	mem(1422) := To_stdlogicvector(X"00");
	mem(1423) := To_stdlogicvector(X"00");
	mem(1424) := To_stdlogicvector(X"00");
	mem(1425) := To_stdlogicvector(X"00");
	mem(1426) := To_stdlogicvector(X"00");
	mem(1427) := To_stdlogicvector(X"00");
	mem(1428) := To_stdlogicvector(X"00");
	mem(1429) := To_stdlogicvector(X"00");
	mem(1430) := To_stdlogicvector(X"00");
	mem(1431) := To_stdlogicvector(X"00");
	mem(1432) := To_stdlogicvector(X"57");
	mem(1433) := To_stdlogicvector(X"E5");
	mem(1434) := To_stdlogicvector(X"00");
	mem(1435) := To_stdlogicvector(X"00");
	mem(1436) := To_stdlogicvector(X"00");
	mem(1437) := To_stdlogicvector(X"00");
	mem(1438) := To_stdlogicvector(X"00");
	mem(1439) := To_stdlogicvector(X"00");
	mem(1440) := To_stdlogicvector(X"00");
	mem(1441) := To_stdlogicvector(X"00");
	mem(1442) := To_stdlogicvector(X"00");
	mem(1443) := To_stdlogicvector(X"00");
	mem(1444) := To_stdlogicvector(X"00");
	mem(1445) := To_stdlogicvector(X"00");
	mem(1446) := To_stdlogicvector(X"80");
	mem(1447) := To_stdlogicvector(X"40");
	mem(1448) := To_stdlogicvector(X"00");
	mem(1449) := To_stdlogicvector(X"00");
	mem(1450) := To_stdlogicvector(X"00");
	mem(1451) := To_stdlogicvector(X"00");
	mem(1452) := To_stdlogicvector(X"00");
	mem(1453) := To_stdlogicvector(X"00");
	mem(1454) := To_stdlogicvector(X"00");
	mem(1455) := To_stdlogicvector(X"00");
	mem(1456) := To_stdlogicvector(X"00");
	mem(1457) := To_stdlogicvector(X"00");
	mem(1458) := To_stdlogicvector(X"00");
	mem(1459) := To_stdlogicvector(X"00");
	mem(1460) := To_stdlogicvector(X"82");
	mem(1461) := To_stdlogicvector(X"73");
	mem(1462) := To_stdlogicvector(X"00");
	mem(1463) := To_stdlogicvector(X"00");
	mem(1464) := To_stdlogicvector(X"00");
	mem(1465) := To_stdlogicvector(X"00");
	mem(1466) := To_stdlogicvector(X"00");
	mem(1467) := To_stdlogicvector(X"00");
	mem(1468) := To_stdlogicvector(X"00");
	mem(1469) := To_stdlogicvector(X"00");
	mem(1470) := To_stdlogicvector(X"00");
	mem(1471) := To_stdlogicvector(X"00");
	mem(1472) := To_stdlogicvector(X"00");
	mem(1473) := To_stdlogicvector(X"00");
	mem(1474) := To_stdlogicvector(X"22");
	mem(1475) := To_stdlogicvector(X"12");
	mem(1476) := To_stdlogicvector(X"00");
	mem(1477) := To_stdlogicvector(X"00");
	mem(1478) := To_stdlogicvector(X"00");
	mem(1479) := To_stdlogicvector(X"00");
	mem(1480) := To_stdlogicvector(X"00");
	mem(1481) := To_stdlogicvector(X"00");
	mem(1482) := To_stdlogicvector(X"00");
	mem(1483) := To_stdlogicvector(X"00");
	mem(1484) := To_stdlogicvector(X"00");
	mem(1485) := To_stdlogicvector(X"00");
	mem(1486) := To_stdlogicvector(X"00");
	mem(1487) := To_stdlogicvector(X"00");
	mem(1488) := To_stdlogicvector(X"A0");
	mem(1489) := To_stdlogicvector(X"5D");
	mem(1490) := To_stdlogicvector(X"00");
	mem(1491) := To_stdlogicvector(X"00");
	mem(1492) := To_stdlogicvector(X"00");
	mem(1493) := To_stdlogicvector(X"00");
	mem(1494) := To_stdlogicvector(X"00");
	mem(1495) := To_stdlogicvector(X"00");
	mem(1496) := To_stdlogicvector(X"00");
	mem(1497) := To_stdlogicvector(X"00");
	mem(1498) := To_stdlogicvector(X"00");
	mem(1499) := To_stdlogicvector(X"00");
	mem(1500) := To_stdlogicvector(X"00");
	mem(1501) := To_stdlogicvector(X"00");
	mem(1502) := To_stdlogicvector(X"0D");
	mem(1503) := To_stdlogicvector(X"04");
	mem(1504) := To_stdlogicvector(X"00");
	mem(1505) := To_stdlogicvector(X"00");
	mem(1506) := To_stdlogicvector(X"00");
	mem(1507) := To_stdlogicvector(X"00");
	mem(1508) := To_stdlogicvector(X"00");
	mem(1509) := To_stdlogicvector(X"00");
	mem(1510) := To_stdlogicvector(X"00");
	mem(1511) := To_stdlogicvector(X"00");
	mem(1512) := To_stdlogicvector(X"00");
	mem(1513) := To_stdlogicvector(X"00");
	mem(1514) := To_stdlogicvector(X"00");
	mem(1515) := To_stdlogicvector(X"00");
	mem(1516) := To_stdlogicvector(X"41");
	mem(1517) := To_stdlogicvector(X"12");
	mem(1518) := To_stdlogicvector(X"00");
	mem(1519) := To_stdlogicvector(X"00");
	mem(1520) := To_stdlogicvector(X"00");
	mem(1521) := To_stdlogicvector(X"00");
	mem(1522) := To_stdlogicvector(X"00");
	mem(1523) := To_stdlogicvector(X"00");
	mem(1524) := To_stdlogicvector(X"00");
	mem(1525) := To_stdlogicvector(X"00");
	mem(1526) := To_stdlogicvector(X"00");
	mem(1527) := To_stdlogicvector(X"00");
	mem(1528) := To_stdlogicvector(X"00");
	mem(1529) := To_stdlogicvector(X"00");
	mem(1530) := To_stdlogicvector(X"0D");
	mem(1531) := To_stdlogicvector(X"ED");
	mem(1532) := To_stdlogicvector(X"00");
	mem(1533) := To_stdlogicvector(X"00");
	mem(1534) := To_stdlogicvector(X"00");
	mem(1535) := To_stdlogicvector(X"00");
	mem(1536) := To_stdlogicvector(X"00");
	mem(1537) := To_stdlogicvector(X"00");
	mem(1538) := To_stdlogicvector(X"00");
	mem(1539) := To_stdlogicvector(X"00");
	mem(1540) := To_stdlogicvector(X"00");
	mem(1541) := To_stdlogicvector(X"00");
	mem(1542) := To_stdlogicvector(X"00");
	mem(1543) := To_stdlogicvector(X"00");
	mem(1544) := To_stdlogicvector(X"83");
	mem(1545) := To_stdlogicvector(X"73");
	mem(1546) := To_stdlogicvector(X"00");
	mem(1547) := To_stdlogicvector(X"00");
	mem(1548) := To_stdlogicvector(X"00");
	mem(1549) := To_stdlogicvector(X"00");
	mem(1550) := To_stdlogicvector(X"00");
	mem(1551) := To_stdlogicvector(X"00");
	mem(1552) := To_stdlogicvector(X"00");
	mem(1553) := To_stdlogicvector(X"00");
	mem(1554) := To_stdlogicvector(X"00");
	mem(1555) := To_stdlogicvector(X"00");
	mem(1556) := To_stdlogicvector(X"00");
	mem(1557) := To_stdlogicvector(X"00");
	mem(1558) := To_stdlogicvector(X"19");
	mem(1559) := To_stdlogicvector(X"E0");
	mem(1560) := To_stdlogicvector(X"00");
	mem(1561) := To_stdlogicvector(X"62");
	mem(1562) := To_stdlogicvector(X"01");
	mem(1563) := To_stdlogicvector(X"64");
	mem(1564) := To_stdlogicvector(X"42");
	mem(1565) := To_stdlogicvector(X"1A");
	mem(1566) := To_stdlogicvector(X"02");
	mem(1567) := To_stdlogicvector(X"7A");
	mem(1568) := To_stdlogicvector(X"03");
	mem(1569) := To_stdlogicvector(X"74");
	mem(1570) := To_stdlogicvector(X"45");
	mem(1571) := To_stdlogicvector(X"1B");
	mem(1572) := To_stdlogicvector(X"82");
	mem(1573) := To_stdlogicvector(X"14");
	mem(1574) := To_stdlogicvector(X"02");
	mem(1575) := To_stdlogicvector(X"7A");
	mem(1576) := To_stdlogicvector(X"03");
	mem(1577) := To_stdlogicvector(X"74");
	mem(1578) := To_stdlogicvector(X"03");
	mem(1579) := To_stdlogicvector(X"6C");
	mem(1580) := To_stdlogicvector(X"02");
	mem(1581) := To_stdlogicvector(X"66");
	mem(1582) := To_stdlogicvector(X"83");
	mem(1583) := To_stdlogicvector(X"17");
	mem(1584) := To_stdlogicvector(X"C3");
	mem(1585) := To_stdlogicvector(X"14");
	mem(1586) := To_stdlogicvector(X"02");
	mem(1587) := To_stdlogicvector(X"52");
	mem(1588) := To_stdlogicvector(X"C2");
	mem(1589) := To_stdlogicvector(X"58");
	mem(1590) := To_stdlogicvector(X"3F");
	mem(1591) := To_stdlogicvector(X"9F");
	mem(1592) := To_stdlogicvector(X"3F");
	mem(1593) := To_stdlogicvector(X"9D");
	mem(1594) := To_stdlogicvector(X"C6");
	mem(1595) := To_stdlogicvector(X"19");
	mem(1596) := To_stdlogicvector(X"FF");
	mem(1597) := To_stdlogicvector(X"0F");
	mem(1598) := To_stdlogicvector(X"00");
	mem(1599) := To_stdlogicvector(X"00");
	mem(1600) := To_stdlogicvector(X"00");
	mem(1601) := To_stdlogicvector(X"00");
	mem(1602) := To_stdlogicvector(X"00");
	mem(1603) := To_stdlogicvector(X"00");
	mem(1604) := To_stdlogicvector(X"00");
	mem(1605) := To_stdlogicvector(X"00");
	mem(1606) := To_stdlogicvector(X"00");
	mem(1607) := To_stdlogicvector(X"00");
	mem(1608) := To_stdlogicvector(X"00");
	mem(1609) := To_stdlogicvector(X"00");
	mem(1610) := To_stdlogicvector(X"09");
	mem(1611) := To_stdlogicvector(X"00");
	mem(1612) := To_stdlogicvector(X"CF");
	mem(1613) := To_stdlogicvector(X"70");
	mem(1614) := To_stdlogicvector(X"00");
	mem(1615) := To_stdlogicvector(X"00");
	mem(1616) := To_stdlogicvector(X"00");
	mem(1617) := To_stdlogicvector(X"00");
	mem(1618) := To_stdlogicvector(X"FF");
	mem(1619) := To_stdlogicvector(X"9D");
	mem(1620) := To_stdlogicvector(X"00");
	mem(1621) := To_stdlogicvector(X"00");
	mem(1622) := To_stdlogicvector(X"00");
	mem(1623) := To_stdlogicvector(X"00");
	mem(1624) := To_stdlogicvector(X"00");
	mem(1625) := To_stdlogicvector(X"00");
	mem(1626) := To_stdlogicvector(X"00");
	mem(1627) := To_stdlogicvector(X"00");
	mem(1628) := To_stdlogicvector(X"00");
	mem(1629) := To_stdlogicvector(X"00");
	mem(1630) := To_stdlogicvector(X"00");
	mem(1631) := To_stdlogicvector(X"00");
	mem(1632) := To_stdlogicvector(X"C0");
	mem(1633) := To_stdlogicvector(X"C1");
	mem(1634) := To_stdlogicvector(X"00");
	mem(1635) := To_stdlogicvector(X"00");
	mem(1636) := To_stdlogicvector(X"00");
	mem(1637) := To_stdlogicvector(X"00");
	mem(1638) := To_stdlogicvector(X"00");
	mem(1639) := To_stdlogicvector(X"00");
	mem(1640) := To_stdlogicvector(X"00");
	mem(1641) := To_stdlogicvector(X"00");
	mem(1642) := To_stdlogicvector(X"00");
	mem(1643) := To_stdlogicvector(X"00");
	mem(1644) := To_stdlogicvector(X"00");
	mem(1645) := To_stdlogicvector(X"00");
	mem(1646) := To_stdlogicvector(X"08");
	mem(1647) := To_stdlogicvector(X"62");
	mem(1648) := To_stdlogicvector(X"00");
	mem(1649) := To_stdlogicvector(X"00");
	mem(1650) := To_stdlogicvector(X"00");
	mem(1651) := To_stdlogicvector(X"00");
	mem(1652) := To_stdlogicvector(X"00");
	mem(1653) := To_stdlogicvector(X"00");
	mem(1654) := To_stdlogicvector(X"00");
	mem(1655) := To_stdlogicvector(X"00");
	mem(1656) := To_stdlogicvector(X"00");
	mem(1657) := To_stdlogicvector(X"00");
	mem(1658) := To_stdlogicvector(X"00");
	mem(1659) := To_stdlogicvector(X"00");
	mem(1660) := To_stdlogicvector(X"06");
	mem(1661) := To_stdlogicvector(X"22");
	mem(1662) := To_stdlogicvector(X"00");
	mem(1663) := To_stdlogicvector(X"00");
	mem(1664) := To_stdlogicvector(X"00");
	mem(1665) := To_stdlogicvector(X"00");
	mem(1666) := To_stdlogicvector(X"00");
	mem(1667) := To_stdlogicvector(X"00");
	mem(1668) := To_stdlogicvector(X"00");
	mem(1669) := To_stdlogicvector(X"00");
	mem(1670) := To_stdlogicvector(X"00");
	mem(1671) := To_stdlogicvector(X"00");
	mem(1672) := To_stdlogicvector(X"00");
	mem(1673) := To_stdlogicvector(X"00");
	mem(1674) := To_stdlogicvector(X"08");
	mem(1675) := To_stdlogicvector(X"24");
	mem(1676) := To_stdlogicvector(X"00");
	mem(1677) := To_stdlogicvector(X"00");
	mem(1678) := To_stdlogicvector(X"00");
	mem(1679) := To_stdlogicvector(X"00");
	mem(1680) := To_stdlogicvector(X"00");
	mem(1681) := To_stdlogicvector(X"00");
	mem(1682) := To_stdlogicvector(X"00");
	mem(1683) := To_stdlogicvector(X"00");
	mem(1684) := To_stdlogicvector(X"00");
	mem(1685) := To_stdlogicvector(X"00");
	mem(1686) := To_stdlogicvector(X"00");
	mem(1687) := To_stdlogicvector(X"00");
	mem(1688) := To_stdlogicvector(X"06");
	mem(1689) := To_stdlogicvector(X"66");
	mem(1690) := To_stdlogicvector(X"00");
	mem(1691) := To_stdlogicvector(X"00");
	mem(1692) := To_stdlogicvector(X"00");
	mem(1693) := To_stdlogicvector(X"00");
	mem(1694) := To_stdlogicvector(X"00");
	mem(1695) := To_stdlogicvector(X"00");
	mem(1696) := To_stdlogicvector(X"00");
	mem(1697) := To_stdlogicvector(X"00");
	mem(1698) := To_stdlogicvector(X"00");
	mem(1699) := To_stdlogicvector(X"00");
	mem(1700) := To_stdlogicvector(X"00");
	mem(1701) := To_stdlogicvector(X"00");
	mem(1702) := To_stdlogicvector(X"00");
	mem(1703) := To_stdlogicvector(X"68");
	mem(1704) := To_stdlogicvector(X"00");
	mem(1705) := To_stdlogicvector(X"00");
	mem(1706) := To_stdlogicvector(X"00");
	mem(1707) := To_stdlogicvector(X"00");
	mem(1708) := To_stdlogicvector(X"00");
	mem(1709) := To_stdlogicvector(X"00");
	mem(1710) := To_stdlogicvector(X"00");
	mem(1711) := To_stdlogicvector(X"00");
	mem(1712) := To_stdlogicvector(X"00");
	mem(1713) := To_stdlogicvector(X"00");
	mem(1714) := To_stdlogicvector(X"00");
	mem(1715) := To_stdlogicvector(X"00");
