	mem(0) := To_stdlogicvector(X"2F");
	mem(1) := To_stdlogicvector(X"19");
	mem(2) := To_stdlogicvector(X"67");
	mem(3) := To_stdlogicvector(X"1B");
	mem(4) := To_stdlogicvector(X"AB");
	mem(5) := To_stdlogicvector(X"1D");
	mem(6) := To_stdlogicvector(X"14");
	mem(7) := To_stdlogicvector(X"62");
	mem(8) := To_stdlogicvector(X"15");
	mem(9) := To_stdlogicvector(X"64");
	mem(10) := To_stdlogicvector(X"16");
	mem(11) := To_stdlogicvector(X"66");
	mem(12) := To_stdlogicvector(X"40");
	mem(13) := To_stdlogicvector(X"6E");
	mem(14) := To_stdlogicvector(X"41");
	mem(15) := To_stdlogicvector(X"7A");
	mem(16) := To_stdlogicvector(X"80");
	mem(17) := To_stdlogicvector(X"6E");
	mem(18) := To_stdlogicvector(X"84");
	mem(19) := To_stdlogicvector(X"7A");
	mem(20) := To_stdlogicvector(X"40");
	mem(21) := To_stdlogicvector(X"6E");
	mem(22) := To_stdlogicvector(X"C1");
	mem(23) := To_stdlogicvector(X"7C");
	mem(24) := To_stdlogicvector(X"81");
	mem(25) := To_stdlogicvector(X"6E");
	mem(26) := To_stdlogicvector(X"C5");
	mem(27) := To_stdlogicvector(X"7C");
	mem(28) := To_stdlogicvector(X"82");
	mem(29) := To_stdlogicvector(X"6E");
	mem(30) := To_stdlogicvector(X"47");
	mem(31) := To_stdlogicvector(X"78");
	mem(32) := To_stdlogicvector(X"84");
	mem(33) := To_stdlogicvector(X"68");
	mem(34) := To_stdlogicvector(X"47");
	mem(35) := To_stdlogicvector(X"68");
	mem(36) := To_stdlogicvector(X"43");
	mem(37) := To_stdlogicvector(X"3A");
	mem(38) := To_stdlogicvector(X"FF");
	mem(39) := To_stdlogicvector(X"0F");
	mem(40) := To_stdlogicvector(X"40");
	mem(41) := To_stdlogicvector(X"00");
	mem(42) := To_stdlogicvector(X"C0");
	mem(43) := To_stdlogicvector(X"00");
	mem(44) := To_stdlogicvector(X"40");
	mem(45) := To_stdlogicvector(X"01");
	mem(46) := To_stdlogicvector(X"00");
	mem(47) := To_stdlogicvector(X"00");
	mem(48) := To_stdlogicvector(X"00");
	mem(49) := To_stdlogicvector(X"00");
	mem(50) := To_stdlogicvector(X"00");
	mem(51) := To_stdlogicvector(X"00");
	mem(64) := To_stdlogicvector(X"11");
	mem(65) := To_stdlogicvector(X"11");
	mem(66) := To_stdlogicvector(X"00");
	mem(67) := To_stdlogicvector(X"00");
	mem(68) := To_stdlogicvector(X"00");
	mem(69) := To_stdlogicvector(X"00");
	mem(70) := To_stdlogicvector(X"00");
	mem(71) := To_stdlogicvector(X"00");
	mem(72) := To_stdlogicvector(X"00");
	mem(73) := To_stdlogicvector(X"00");
	mem(74) := To_stdlogicvector(X"00");
	mem(75) := To_stdlogicvector(X"00");
	mem(76) := To_stdlogicvector(X"00");
	mem(77) := To_stdlogicvector(X"00");
	mem(78) := To_stdlogicvector(X"00");
	mem(79) := To_stdlogicvector(X"00");
	mem(192) := To_stdlogicvector(X"22");
	mem(193) := To_stdlogicvector(X"22");
	mem(194) := To_stdlogicvector(X"00");
	mem(195) := To_stdlogicvector(X"00");
	mem(196) := To_stdlogicvector(X"00");
	mem(197) := To_stdlogicvector(X"00");
	mem(198) := To_stdlogicvector(X"00");
	mem(199) := To_stdlogicvector(X"00");
	mem(200) := To_stdlogicvector(X"00");
	mem(201) := To_stdlogicvector(X"00");
	mem(202) := To_stdlogicvector(X"00");
	mem(203) := To_stdlogicvector(X"00");
	mem(204) := To_stdlogicvector(X"00");
	mem(205) := To_stdlogicvector(X"00");
	mem(206) := To_stdlogicvector(X"00");
	mem(207) := To_stdlogicvector(X"00");
	mem(320) := To_stdlogicvector(X"33");
	mem(321) := To_stdlogicvector(X"33");
	mem(322) := To_stdlogicvector(X"00");
	mem(323) := To_stdlogicvector(X"00");
	mem(324) := To_stdlogicvector(X"00");
	mem(325) := To_stdlogicvector(X"00");
	mem(326) := To_stdlogicvector(X"00");
	mem(327) := To_stdlogicvector(X"00");
	mem(328) := To_stdlogicvector(X"00");
	mem(329) := To_stdlogicvector(X"00");
	mem(330) := To_stdlogicvector(X"00");
	mem(331) := To_stdlogicvector(X"00");
	mem(332) := To_stdlogicvector(X"00");
	mem(333) := To_stdlogicvector(X"00");
	mem(334) := To_stdlogicvector(X"00");
	mem(335) := To_stdlogicvector(X"00");
